netcdf \2014-12-04 {
dimensions:
	ts_dim = 1 ;
	layer_dim = 23062 ;
	descriptChar = 214 ;
	familyidChar = 33 ;
	site_noChar = 15 ;
	station_nmChar = 50 ;
	site_tp_cdChar = 6 ;
	dec_coord_datum_cdChar = 5 ;
	alt_datum_cdChar = 7 ;
	huc_cdChar = 8 ;
	tz_cdChar = 4 ;
	agency_cdChar = 5 ;
	district_cdChar = 3 ;
	county_cdChar = 3 ;
	country_cdChar = 2 ;
variables:
	int time(ts_dim) ;
	double v00060_value(ts_dim, layer_dim) ;
	double v00065_value(ts_dim, layer_dim) ;
	double v00010_value(ts_dim, layer_dim) ;
	double v00095_value(ts_dim, layer_dim) ;
	double v00035_value(ts_dim, layer_dim) ;
	double v00036_value(ts_dim, layer_dim) ;
	double v00045_value(ts_dim, layer_dim) ;
	double v00062_value(ts_dim, layer_dim) ;
	double v00054_value(ts_dim, layer_dim) ;
	double v00060_validated(ts_dim, layer_dim) ;
	double v00065_validated(ts_dim, layer_dim) ;
	double v00010_validated(ts_dim, layer_dim) ;
	double v00095_validated(ts_dim, layer_dim) ;
	double v00035_validated(ts_dim, layer_dim) ;
	double v00036_validated(ts_dim, layer_dim) ;
	double v00045_validated(ts_dim, layer_dim) ;
	double v00062_validated(ts_dim, layer_dim) ;
	double v00054_validated(ts_dim, layer_dim) ;
	char v00060_description(layer_dim, descriptChar) ;
	char v00065_description(layer_dim, descriptChar) ;
	char v00010_description(layer_dim, descriptChar) ;
	char v00095_description(layer_dim, descriptChar) ;
	char v00035_description(layer_dim, descriptChar) ;
	char v00036_description(layer_dim, descriptChar) ;
	char v00045_description(layer_dim, descriptChar) ;
	char v00062_description(layer_dim, descriptChar) ;
	char v00054_description(layer_dim, descriptChar) ;
	char familyid(layer_dim, familyidChar) ;
	char site_no(layer_dim, site_noChar) ;
	int dd_nu(layer_dim) ;
	char station_nm(layer_dim, station_nmChar) ;
	char site_tp_cd(layer_dim, site_tp_cdChar) ;
	double dec_lat_va(layer_dim) ;
	double dec_long_va(layer_dim) ;
	char dec_coord_datum_cd(layer_dim, dec_coord_datum_cdChar) ;
	double alt_va(layer_dim) ;
	char alt_datum_cd(layer_dim, alt_datum_cdChar) ;
	char huc_cd(layer_dim, huc_cdChar) ;
	char tz_cd(layer_dim, tz_cdChar) ;
	char agency_cd(layer_dim, agency_cdChar) ;
	char district_cd(layer_dim, district_cdChar) ;
	char county_cd(layer_dim, county_cdChar) ;
	char country_cd(layer_dim, country_cdChar) ;
data:

 time = 1417651200 ;

 v00060_value =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 288, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 288, 1, 96, 1, 
    1, 288, 1, 85, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 288, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 288, 96, 1, 96, 1, 96, 1, 96, 1, 1, 86, 1, 92, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 95, 1, 1, 1, 96, 96, 1, 1, 96, 96, 
    1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 132, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 93, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 89, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 
    1, 144, 1, 1, 1, 151, 1, 1, 1, 87, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 144, 
    1, 1, 1, 111, 1, 1, 1, 144, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 73, 1, 96, 1, 1, 96, 96, 1, 95, 
    1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 144, 1, 144, 1, 1, 1, 1, 1, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 144, 1, 144, 1, 1, 1, 1, 1, 144, 1, 144, 1, 1, 1, 
    1, 1, 144, 1, 1, 1, 144, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    144, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 95, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 288, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 95, 1, 1, 96, 84, 1, 96, 1, 96, 1, 1, 96, 1, 95, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 95, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 91, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 1, 288, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 94, 1, 1, 1, 
    1, 96, 1, 1, 96, 96, 1, 288, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    288, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 288, 1, 96, 1, 96, 96, 1, 1, 1, 288, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 95, 96, 1, 96, 1, 1, 1, 96, 1, 288, 1, 96, 1, 96, 96, 1, 1, 1, 96, 
    1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 240, 1, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 288, 96, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 288, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 52, 1, 
    1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 288, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 95, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 288, 1, 1, 1, 1, 1, 40, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 288, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 288, 1, 96, 1, 288, 1, 288, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 288, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 240, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 240, 1, 96, 1, 1, 240, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 
    288, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 95, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 96, 1, 
    1, 48, 1, 1, 1, 96, 96, 1, 1, 1, 1, 48, 1, 1, 96, 1, 48, 1, 1, 1, 96, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 288, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 96, 1, 1, 96, 96, 1, 1, 92, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 53, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 240, 1, 1, 240, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 95, 1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 
    92, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 48, 1, 96, 96, 1, 1, 1, 1, 48, 1, 96, 1, 96, 1, 1, 48, 1, 1, 
    96, 48, 1, 1, 1, 1, 96, 1, 94, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 95, 95, 1, 
    1, 1, 96, 1, 96, 1, 1, 48, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 
    96, 96, 1, 1, 288, 1, 1, 1, 1, 1, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 288, 1, 1, 288, 1, 
    243, 96, 1, 96, 1, 1, 288, 96, 1, 1, 96, 288, 1, 1, 288, 1, 1439, 1, 
    1440, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 288, 1, 1, 96, 1, 
    96, 1, 96, 1, 288, 96, 1, 1, 288, 1, 166, 1, 1, 288, 1, 288, 1, 288, 288, 
    1, 1, 288, 96, 1, 1, 720, 96, 1, 1, 288, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 288, 1, 288, 96, 1, 96, 1, 95, 1, 96, 1, 1, 96, 1, 96, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 92, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 94, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 
    288, 96, 1, 96, 1, 95, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 288, 1, 288, 
    1, 288, 1, 288, 1, 288, 1, 96, 96, 1, 1, 288, 1, 1, 1, 288, 1, 1, 96, 1, 
    1, 1, 1, 288, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 288, 1, 288, 1, 
    1, 288, 1, 1, 1, 96, 1, 1, 288, 1, 1, 96, 1, 1, 288, 1, 288, 1, 96, 1, 1, 
    288, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 288, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 288, 1, 1, 96, 1, 1, 
    288, 1, 1, 95, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 288, 1, 1, 96, 288, 1, 1, 
    1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 95, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 66, 1, 1, 1, 1, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 288, 1, 288, 1, 288, 1, 96, 1, 288, 1, 1, 288, 1, 288, 1, 96, 1, 
    288, 1, 288, 1, 288, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 48, 1, 1, 48, 1, 1, 96, 24, 1, 1, 1, 96, 96, 1, 
    1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 288, 1, 288, 1, 288, 1, 288, 1, 
    96, 288, 1, 1, 288, 1, 288, 1, 288, 1, 288, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 288, 1, 1, 288, 1, 288, 288, 1, 1, 
    288, 1, 1, 288, 1, 288, 1, 1, 288, 1, 1, 288, 1, 1, 288, 1, 1, 1, 288, 1, 
    288, 1, 288, 288, 1, 288, 1, 1, 288, 1, 288, 1, 288, 1, 288, 288, 1, 1, 
    1, 1, 288, 1, 288, 1, 1, 288, 1, 288, 1, 96, 1, 288, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 24, 1, 1, 96, 1, 96, 1, 96, 1, 1, 24, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 96, 1, 96, 1, 96, 24, 
    1, 1, 1, 24, 96, 1, 1, 24, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 91, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 24, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 72, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 95, 1, 1, 95, 1, 96, 1, 1, 95, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 94, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 94, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 24, 
    96, 1, 96, 1, 1, 48, 24, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 1, 1, 1, 95, 94, 1, 1, 96, 96, 1, 96, 1, 1, 83, 1, 1, 96, 1, 
    48, 1, 48, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 48, 1, 24, 1, 24, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 24, 1, 1, 1, 1, 48, 96, 1, 1, 1, 24, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    24, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    24, 1, 48, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 288, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 48, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 24, 1, 1, 48, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 221, 1, 1, 96, 1, 89, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 264, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 
    1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 95, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 84, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 96, 24, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 96, 1, 1, 1, 1, 1, 87, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 203, 1, 1, 1, 1, 1, 1, 1, 24, 1, 24, 1, 24, 1, 92, 1, 24, 
    1, 24, 1, 1, 95, 96, 1, 1, 96, 96, 1, 96, 1, 1, 24, 48, 1, 48, 1, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 24, 1, 24, 1, 1, 24, 1, 
    96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 
    92, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 24, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 24, 1, 1, 24, 24, 1, 1, 1, 1, 24, 1, 96, 1, 24, 1, 96, 1, 1, 
    96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 24, 1, 1, 24, 1, 23, 1, 24, 1, 
    1, 24, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 24, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 24, 1, 1, 24, 1, 24, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 91, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 95, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 92, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 93, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 24, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 94, 1, 1, 92, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 48, 24, 
    1, 1, 96, 1, 1, 48, 48, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 48, 1, 24, 1, 1, 
    96, 1, 1, 1, 24, 1, 1, 48, 24, 1, 1, 48, 48, 1, 96, 1, 1, 96, 1, 96, 48, 
    1, 48, 1, 96, 1, 48, 1, 96, 1, 1, 96, 1, 48, 1, 48, 1, 96, 1, 24, 1, 48, 
    1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 48, 1, 1, 48, 1, 48, 96, 1, 96, 
    1, 1, 1, 48, 1, 48, 1, 96, 1, 24, 1, 1, 48, 1, 1, 96, 1, 48, 48, 1, 1, 
    96, 1, 1, 56, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 95, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 95, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 48, 1, 48, 1, 1, 48, 
    1, 1, 1, 1, 96, 48, 1, 48, 1, 1, 48, 1, 48, 1, 48, 1, 1, 48, 1, 1, 96, 
    96, 1, 1, 96, 1, 1, 1, 48, 1, 1, 1, 48, 48, 1, 95, 1, 1, 1, 96, 1, 48, 1, 
    48, 1, 48, 1, 47, 1, 1, 96, 1, 96, 24, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 
    48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 44, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 24, 1, 1, 48, 
    1, 1, 24, 1, 1, 1, 1, 96, 24, 1, 1, 1, 96, 1, 96, 1, 96, 1, 24, 1, 1, 96, 
    96, 1, 1, 1, 96, 1, 80, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 24, 1, 1, 24, 
    1, 96, 1, 1, 1, 96, 24, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 48, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 288, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 96, 1, 96, 1, 1, 90, 1, 1, 48, 1, 1, 24, 1, 1, 48, 1, 1, 1, 48, 1, 
    96, 1, 48, 1, 96, 1, 48, 1, 93, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 25, 1, 96, 1, 93, 1, 1, 1, 95, 1, 96, 1, 82, 1, 96, 1, 1, 81, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 24, 1, 1, 48, 1, 48, 1, 48, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 91, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 95, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 89, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    24, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 48, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 48, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 93, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 48, 1, 1, 95, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 95, 1, 1, 96, 1, 95, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 84, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 288, 1, 96, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 48, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 24, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 
    1, 1, 95, 1, 1, 1, 1, 96, 96, 1, 1, 48, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 1, 1, 48, 1, 48, 1, 96, 1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 96, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 96, 
    1, 1, 48, 1, 1, 1, 96, 1, 48, 1, 1, 24, 48, 1, 1, 96, 1, 1, 1, 48, 1, 96, 
    1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 96, 1, 1, 48, 1, 63, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 96, 1, 1, 96, 1, 1, 1, 48, 1, 
    96, 1, 1, 1, 96, 1, 48, 1, 48, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 48, 
    1, 1, 48, 1, 1, 96, 1, 1, 96, 1, 1, 1, 48, 1, 1, 96, 1, 48, 1, 1, 96, 1, 
    1, 95, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 48, 48, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 48, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 48, 1, 1, 1, 1, 46, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 1, 42, 1, 1, 
    1, 48, 1, 1, 47, 1, 1, 1, 47, 1, 1, 1, 96, 1, 48, 1, 48, 48, 1, 1, 1, 1, 
    96, 1, 1, 1, 48, 1, 48, 1, 48, 1, 1, 1, 48, 1, 48, 1, 96, 1, 48, 1, 1, 
    96, 1, 48, 48, 1, 1, 48, 1, 1, 1, 48, 1, 47, 1, 1, 1, 1, 48, 46, 1, 1, 
    96, 1, 48, 24, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 48, 1, 1, 1, 96, 96, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 
    1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 288, 1, 1, 288, 1, 1, 264, 1, 1, 96, 1, 
    1, 95, 1, 1, 92, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 288, 1, 1, 
    288, 1, 1, 96, 1, 96, 1, 288, 1, 1, 288, 288, 1, 1, 1, 288, 1, 1, 1, 288, 
    1, 288, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 144, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 93, 1, 1, 1, 96, 1, 1, 92, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    95, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 92, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 1, 90, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 95, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 95, 96, 1, 1, 1, 1, 1, 1, 1, 48, 1, 
    48, 1, 1, 1, 48, 96, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 48, 1, 1, 
    1, 48, 1, 1, 48, 92, 1, 96, 1, 1, 1, 48, 1, 1, 1, 96, 1, 1, 1, 96, 48, 1, 
    1, 1, 1, 1, 48, 1, 1, 91, 1, 48, 1, 1, 1, 1, 1, 48, 1, 48, 1, 1, 1, 48, 
    48, 1, 1, 1, 1, 1, 97, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 97, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 94, 1, 1, 1, 1, 
    1, 1, 97, 1, 1, 97, 1, 1, 96, 1, 48, 1, 96, 1, 1, 96, 96, 1, 1, 48, 1, 1, 
    43, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 48, 1, 1, 1, 1, 48, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 48, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 48, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 48, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 48, 1, 95, 1, 1, 96, 1, 96, 
    96, 1, 48, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 
    1, 1, 48, 1, 96, 1, 1, 96, 1, 48, 1, 1, 1, 96, 96, 1, 1, 95, 1, 1, 288, 
    1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 93, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 24, 1, 1, 96, 96, 1, 1, 22, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 24, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 
    96, 1, 1, 94, 1, 96, 1, 96, 1, 1, 96, 1, 1, 24, 1, 96, 24, 1, 1, 96, 1, 
    96, 96, 1, 1, 1, 96, 1, 24, 49, 1, 1, 96, 1, 96, 1, 1, 1, 1, 48, 1, 1, 
    288, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 9, 1, 1, 1, 96, 1, 288, 
    1, 288, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 24, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 288, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 288, 1, 1, 96, 1, 1, 288, 1, 1, 1, 96, 1, 135, 1, 96, 
    1, 1, 1, 288, 1, 1, 96, 1, 1, 34, 1, 1, 95, 1, 1, 96, 1, 1, 288, 96, 1, 
    96, 1, 1, 1, 93, 1, 1, 1, 96, 1, 1, 288, 1, 1, 1, 288, 1, 1, 96, 1, 1, 1, 
    1, 288, 1, 1, 288, 1, 1, 288, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 264, 287, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 288, 1, 1, 96, 1, 1, 273, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 48, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 120, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 92, 1, 96, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 120, 
    1, 1, 1, 120, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 45, 1, 1, 240, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 288, 96, 1, 1, 96, 96, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 48, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 
    96, 1, 1, 48, 1, 1, 48, 1, 97, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 48, 96, 1, 1, 96, 1, 
    93, 1, 1, 48, 1, 48, 1, 1, 48, 1, 48, 48, 1, 96, 1, 1, 48, 1, 96, 96, 1, 
    1, 1, 48, 1, 96, 1, 96, 1, 48, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 288, 1, 
    1, 96, 1, 48, 1, 96, 1, 96, 1, 96, 1, 288, 1, 96, 1, 96, 1, 288, 96, 1, 
    1, 1, 1, 48, 1, 1, 96, 1, 1, 144, 1, 96, 1, 1, 1, 48, 1, 48, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 99, 1, 99, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 97, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 98, 1, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 1, 288, 1, 288, 96, 1, 94, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 81, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 26, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 10, 1, 
    96, 1, 95, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 89, 1, 1, 96, 
    1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 48, 1, 48, 1, 96, 1, 96, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 74, 1, 96, 1, 96, 1, 48, 96, 
    1, 48, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 25, 1, 1, 1, 96, 1, 88, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 47, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 82, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 14, 1, 1, 96, 1, 
    24, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 95, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    288, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 88, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 87, 57, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 144, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    288, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 288, 1, 96, 96, 1, 96, 1, 96, 1, 
    288, 1, 1, 1, 288, 96, 1, 1, 1, 1, 1, 288, 1, 96, 1, 1, 1, 288, 1, 1, 96, 
    1, 1, 1, 1, 189, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 144, 
    1, 1, 1, 96, 1, 1, 1, 288, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 90, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 81, 1, 96, 1, 96, 1, 96, 1, 1, 82, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 86, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 13, 90, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 92, 1, 96, 1, 1, 1, 96, 96, 1, 1, 8, 96, 1, 
    96, 1, 96, 1, 144, 1, 96, 1, 58, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 48, 48, 1, 1, 96, 1, 1, 47, 
    46, 1, 1, 1, 48, 1, 48, 1, 48, 1, 48, 1, 48, 1, 1, 1, 1, 48, 1, 1, 48, 
    96, 1, 48, 1, 1, 1, 288, 1, 1, 288, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 95, 1, 95, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 1, 96, 96, 1, 95, 1, 1, 1, 288, 1, 1, 1, 96, 1, 1, 288, 1, 1, 1, 
    1, 288, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 95, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 144, 1, 144, 1, 1, 1, 96, 1, 48, 1, 1, 96, 1, 1, 288, 1, 
    278, 1, 1, 96, 1, 96, 1, 1, 288, 1, 288, 1, 288, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 288, 1, 96, 
    1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 288, 1, 288, 1, 1, 
    1, 75, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 24, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 286, 1, 1, 96, 1, 1, 96, 96, 1, 1, 93, 1, 
    96, 1, 96, 1, 94, 48, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 95, 1, 96, 1, 96, 95, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 94, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 
    1, 1, 69, 1, 49, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 58, 
    96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 95, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 61, 1, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 34, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 35, 1, 1, 86, 1, 96, 
    1, 1, 96, 96, 1, 96, 1, 95, 1, 96, 1, 1, 88, 1, 96, 96, 1, 1, 96, 1, 96, 
    94, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 50, 1, 1, 96, 96, 1, 
    96, 1, 73, 1, 1, 96, 57, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 95, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 37, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 95, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 92, 1, 84, 1, 32, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 288, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 288, 1, 1, 288, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 88, 1, 96, 1, 96, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 288, 1, 288, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 95, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 62, 
    1, 96, 89, 1, 96, 1, 1, 96, 1, 1, 1, 1, 92, 1, 96, 1, 1, 1, 1, 96, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 87, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 95, 1, 1, 1, 
    1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 70, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 14, 1, 1, 1, 96, 1, 96, 1, 1, 49, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 25, 1, 1, 96, 
    1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 33, 1, 1, 97, 1, 
    1, 1, 1, 1, 1, 93, 1, 1, 1, 1, 89, 1, 1, 88, 1, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 88, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 
    1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 96, 1, 288, 1, 1, 288, 1, 288, 96, 
    1, 1, 1, 288, 1, 288, 1, 1, 288, 1, 288, 1, 288, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 288, 1, 42, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 288, 
    1, 288, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 288, 1, 1, 172, 1, 96, 96, 1, 
    1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    29, 1, 1, 94, 96, 1, 1, 89, 96, 1, 1, 96, 95, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 95, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 90, 1, 96, 1, 1, 71, 1, 
    95, 96, 1, 1, 1, 96, 1, 96, 1, 52, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 
    1, 49, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 288, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 
    1, 96, 1, 94, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 95, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 81, 1, 96, 96, 1, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 88, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 90, 1, 1, 
    288, 1, 1, 4, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 94, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 89, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 92, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 69, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 54, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 36, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 94, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 97, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 94, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 288, 1, 288, 1, 1, 288, 
    1, 264, 92, 1, 1, 1, 288, 96, 1, 1, 1, 288, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 288, 1, 1, 288, 1, 288, 288, 1, 1, 1, 288, 1, 
    288, 1, 24, 1, 1, 1, 1, 1, 281, 1, 288, 288, 1, 1, 1, 287, 1, 288, 1, 
    288, 1, 288, 1, 1, 24, 288, 1, 1, 285, 1, 288, 1, 1, 264, 1, 288, 1, 288, 
    1, 288, 288, 1, 1, 288, 1, 1, 264, 1, 290, 288, 1, 1, 288, 288, 1, 1, 96, 
    1, 1, 1, 48, 1, 96, 1, 1, 1, 48, 96, 1, 1, 1, 47, 1, 96, 1, 1, 1, 48, 94, 
    1, 1, 1, 48, 264, 1, 1, 288, 1, 1, 1, 288, 1, 288, 288, 1, 1, 1, 288, 
    255, 1, 1, 287, 1, 48, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 46, 1, 96, 1, 1, 
    94, 96, 1, 24, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 48, 
    1, 1, 24, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 1, 48, 1, 24, 1, 48, 1, 1, 1, 24, 
    96, 1, 1, 1, 1, 277, 89, 1, 24, 1, 1, 1, 288, 1, 1, 288, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 288, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    22, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 95, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 98, 1, 1, 96, 
    47, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 92, 1, 1, 55, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 
    1, 1, 1, 96, 24, 1, 1, 96, 1, 1, 1, 24, 1, 1, 286, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 156, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 85, 1, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 86, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 
    1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 48, 1, 1, 96, 1, 48, 1, 1, 24, 48, 1, 1, 1, 96, 1, 
    1, 1, 48, 1, 96, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 96, 48, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 24, 1, 1, 48, 1, 1, 96, 1, 92, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 24, 1, 1, 1, 96, 1, 96, 96, 
    1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 48, 1, 96, 1, 1, 48, 1, 1, 96, 1, 1, 26, 
    1, 1, 1, 1, 96, 1, 96, 1, 48, 1, 48, 1, 1, 1, 1, 1, 48, 24, 1, 1, 95, 1, 
    96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 70, 1, 48, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 48, 1, 1, 24, 1, 1, 1, 
    96, 92, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 94, 1, 96, 1, 1, 
    24, 96, 1, 48, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 48, 1, 1, 96, 1, 1, 94, 1, 1, 48, 1, 1, 96, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 96, 
    1, 1, 1, 288, 1, 96, 1, 1, 1, 1, 290, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 24, 1, 96, 1, 1, 96, 1, 1, 96, 1, 48, 1, 1, 96, 1, 1, 24, 1, 1, 
    96, 1, 48, 1, 1, 96, 1, 1, 1, 1, 1, 48, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 92, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 48, 1, 1, 48, 48, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 1, 96, 48, 1, 1, 1, 1, 48, 96, 1, 
    1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 24, 
    1, 48, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 
    48, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 48, 1, 1, 1, 
    48, 1, 96, 1, 1, 48, 1, 1, 1, 96, 1, 48, 1, 48, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 93, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 70, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 1, 1, 
    30, 1, 24, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    15, 1, 1, 96, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 86, 1, 1, 60, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 
    1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    96, 1, 48, 1, 1, 48, 1, 1, 1, 48, 1, 48, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    62, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 93, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 48, 1, 37, 1, 1, 1, 48, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 48, 1, 48, 1, 1, 96, 1, 1, 95, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 48, 1, 1, 96, 1, 96, 1, 96, 48, 1, 1, 1, 96, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 144, 1, 24, 1, 1, 1, 1, 96, 24, 1, 1, 1, 
    48, 1, 1, 1, 96, 1, 1, 48, 1, 24, 1, 96, 1, 1, 46, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 24, 96, 96, 1, 1, 1, 1, 24, 1, 
    1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 24, 1, 1, 48, 1, 24, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 90, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 48, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 285, 1, 1, 1, 288, 1, 288, 1, 1, 96, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 24, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 95, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 96, 48, 1, 1, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 48, 1, 1, 48, 1, 1, 48, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 48, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 56, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 48, 1, 1, 48, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 
    1, 1, 1, 1, 1, 40, 48, 1, 1, 48, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 48, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 96, 1, 1, 95, 96, 1, 1, 96, 1, 85, 1, 1, 1, 48, 1, 96, 
    1, 1, 1, 1, 92, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 88, 96, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 95, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 73, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    94, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 94, 96, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 95, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 95, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 87, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 6, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 26, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 60, 1, 1, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 90, 1, 1, 96, 1, 96, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 95, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 95, 1, 1, 288, 1, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 288, 1, 1, 95, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    288, 1, 96, 1, 1, 1, 96, 1, 288, 1, 1, 1, 288, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 288, 1, 1, 288, 95, 
    1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 95, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 288, 
    1, 288, 1, 1, 1, 96, 1, 1, 288, 1, 1, 288, 1, 1, 96, 1, 1, 1, 288, 1, 1, 
    288, 1, 1, 96, 1, 288, 1, 288, 1, 288, 1, 288, 1, 288, 1, 288, 1, 288, 1, 
    288, 1, 1, 288, 96, 1, 1, 1, 1, 288, 1, 288, 288, 1, 1, 288, 1, 288, 288, 
    1, 1, 288, 1, 288, 1, 1, 1, 1, 1, 288, 1, 288, 1, 288, 1, 1, 1, 288, 196, 
    1, 1, 288, 288, 1, 1, 288, 288, 1, 1, 288, 288, 1, 288, 1, 288, 1, 288, 
    1, 288, 1, 1, 288, 1, 1, 96, 288, 1, 1, 1, 288, 1, 1, 1, 1, 96, 1, 1, 96, 
    96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 93, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 95, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 68, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 92, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 95, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 11, 
    1, 1, 96, 288, 1, 1, 1, 96, 1, 1, 96, 96, 1, 288, 1, 288, 1, 1, 1, 96, 1, 
    96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 93, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 
    16, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 144, 1, 
    1, 1, 288, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 95, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 96, 64, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 80, 
    96, 1, 1, 4, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 1, 93, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 93, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 288, 1, 1, 96, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 
    96, 1, 1, 96, 94, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 92, 1, 1, 94, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 90, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 91, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 94, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 101, 1, 1, 1, 
    93, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 94, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 96, 1, 1, 94, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 
    1, 1, 1, 96, 96, 1, 96, 1, 95, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 95, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 192, 
    1, 1, 96, 1, 192, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 81, 1, 96, 1, 
    44, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 65, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 53, 1, 1, 1, 1, 96, 1, 95, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 98, 1, 96, 1, 1, 96, 1, 1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 95, 1, 1, 1, 1, 164, 1, 96, 1, 96, 1, 96, 97, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 100, 1, 96, 96, 1, 99, 1, 96, 1, 1, 96, 96, 1, 1, 97, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 97, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    94, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 62, 96, 1, 1, 96, 96, 96, 96, 96, 96, 
    96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 94, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 92, 1, 90, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 92, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 35, 1, 1, 1, 1, 
    43, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 76, 1, 1, 1, 1, 1, 96, 96, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 80, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 15, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 95, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 89, 1, 96, 1, 76, 1, 96, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 85, 1, 96, 1, 96, 1, 96, 1, 62, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 90, 1, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 95, 1, 96, 1, 1, 95, 1, 1, 1, 98, 1, 96, 
    1, 100, 1, 96, 1, 96, 1, 96, 1, 1, 96, 98, 1, 1, 96, 1, 96, 96, 1, 96, 1, 
    96, 1, 94, 1, 32, 1, 288, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 
    1, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 93, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 49, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 96, 1, 96, 1, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    94, 1, 1, 95, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 85, 1, 85, 1, 85, 1, 85, 1, 1, 85, 86, 1, 
    82, 82, 1, 82, 1, 1, 82, 82, 1, 1, 1, 82, 1, 82, 1, 82, 1, 86, 1, 96, 1, 
    96, 1, 1, 96, 86, 1, 86, 1, 86, 1, 86, 87, 1, 59, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 93, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 84, 1, 1, 1, 84, 1, 84, 1, 78, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 96, 96, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 35, 
    1, 1, 96, 1, 96, 1, 1, 1, 84, 1, 84, 1, 1, 1, 1, 84, 84, 1, 1, 1, 84, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 84, 1, 1, 89, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 54, 1, 1, 96, 1, 96, 1, 83, 1, 1, 
    1, 75, 1, 1, 1, 1, 96, 1, 96, 1, 1, 72, 96, 1, 1, 1, 96, 96, 1, 1, 20, 
    96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    60, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 144, 1, 48, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 227, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 144, 1, 144, 1, 144, 1, 144, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 91, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 53, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 32, 1, 86, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 24, 1, 96, 1, 24, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 48, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 95, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 94, 1, 96, 1, 
    66, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 93, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 56, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 288, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 97, 
    1, 96, 95, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 19, 1, 1, 
    96, 1, 96, 1, 96, 1, 43, 1, 11, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 83, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 89, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 97, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 56, 1, 1, 84, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 99, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 41, 1, 96, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 52, 1, 96, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 28, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 44, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 86, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 48, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 89, 1, 
    1, 1, 48, 1, 1, 48, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 98, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 97, 1, 1, 96, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 114, 1, 1, 108, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    106, 1, 96, 1, 1, 1, 96, 1, 1, 112, 1, 1, 1, 1, 107, 1, 1, 1, 1, 1, 1, 1, 
    137, 1, 1, 126, 1, 128, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 94, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 288, 1, 1, 97, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 95, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 1, 48, 1, 96, 1, 1, 42, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 87, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 88, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 15, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 64, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 94, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 225, 96, 1, 96, 1, 96, 1, 96, 1, 
    112, 1, 96, 1, 102, 1, 100, 1, 96, 1, 96, 1, 288, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 52, 96, 1, 1, 1, 1, 14, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 84, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 58, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 137, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 88, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 288, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 890, 1, 1, 96, 1, 1, 96, 1, 89, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 288, 1, 1193, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 88, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1 ;

 v00065_value =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 96, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 288, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 288, 1, 1, 1, 96, 
    288, 1, 85, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 96, 1, 
    96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 288, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 288, 1, 1, 96, 1, 96, 1, 96, 1, 96, 86, 1, 92, 
    1, 1, 96, 1, 96, 96, 1, 92, 96, 1, 96, 1, 1, 95, 96, 96, 1, 1, 96, 96, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 144, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 93, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 89, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 96, 1, 1, 96, 
    1, 96, 144, 1, 1, 1, 151, 1, 1, 1, 87, 1, 1, 1, 97, 1, 1, 1, 1, 1, 1, 1, 
    144, 1, 1, 1, 111, 1, 1, 1, 144, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 73, 1, 96, 96, 1, 
    1, 96, 1, 95, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 
    144, 1, 1, 96, 1, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 144, 
    1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 144, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 95, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 95, 96, 1, 1, 84, 1, 96, 1, 96, 96, 1, 95, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 91, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 288, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 288, 1, 1, 
    1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 94, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 288, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 288, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 96, 1, 96, 1, 96, 96, 1, 48, 45, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 96, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    72, 1, 96, 96, 1, 1, 96, 96, 1, 96, 96, 96, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 96, 1, 288, 1, 96, 1, 96, 1, 1, 96, 
    96, 288, 1, 12, 1, 96, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 
    288, 288, 1, 288, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 95, 1, 1, 96, 1, 
    96, 1, 96, 1, 288, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 96, 1, 1, 96, 240, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 288, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 288, 96, 1, 96, 1, 1, 96, 1, 96, 96, 52, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 288, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 95, 1, 96, 1, 96, 1, 96, 96, 
    96, 1, 96, 1, 1, 288, 1, 1, 288, 1, 1, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 96, 288, 1, 288, 288, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 288, 1, 288, 240, 1, 1, 288, 288, 1, 96, 1, 96, 1, 96, 96, 1, 
    1, 96, 96, 96, 1, 1, 288, 1, 96, 1, 288, 1, 288, 1, 1, 96, 1, 96, 96, 1, 
    96, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 96, 96, 1, 96, 96, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 288, 
    96, 1, 96, 1, 96, 96, 96, 96, 1, 96, 1, 1, 96, 96, 1, 119, 1, 240, 1, 1, 
    96, 1, 96, 185, 1, 1, 96, 1, 96, 240, 1, 1, 96, 96, 1, 1, 1, 240, 1, 1, 
    96, 240, 1, 240, 1, 1, 1, 96, 96, 1, 240, 1, 1, 240, 1, 1, 1, 96, 240, 1, 
    1, 240, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 240, 1, 240, 1, 230, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 96, 240, 1, 240, 1, 237, 1, 240, 1, 240, 1, 
    240, 1, 240, 1, 96, 1, 1, 96, 240, 1, 96, 206, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 
    1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 288, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 
    96, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 96, 96, 1, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 95, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 1, 
    96, 1, 1, 48, 1, 96, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 96, 1, 48, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 288, 1, 96, 96, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 92, 1, 240, 1, 1, 239, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 53, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 240, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 96, 240, 1, 1, 1, 1, 1, 1, 240, 1, 96, 1, 96, 1, 1, 240, 240, 1, 
    1, 240, 96, 1, 240, 240, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 
    240, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 
    1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 95, 
    1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 
    1, 96, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 96, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 92, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 48, 1, 96, 1, 1, 96, 1, 1, 
    48, 1, 96, 1, 96, 1, 1, 48, 1, 1, 96, 1, 1, 48, 1, 1, 96, 1, 94, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 95, 1, 1, 95, 1, 1, 1, 96, 1, 96, 48, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    1, 1, 96, 96, 1, 240, 240, 96, 1, 1, 96, 96, 1, 1, 96, 288, 1, 1, 1, 1, 
    1, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 288, 288, 1, 243, 1, 1, 96, 1, 96, 288, 1, 1, 
    96, 96, 1, 1, 288, 288, 1, 1439, 1, 1440, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 96, 1, 1, 288, 96, 1, 96, 1, 96, 1, 288, 1, 1, 96, 288, 1, 
    166, 1, 288, 288, 1, 288, 1, 288, 1, 1, 288, 288, 1, 1, 96, 720, 1, 1, 
    96, 288, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 288, 1, 288, 1, 1, 96, 
    1, 96, 1, 95, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 288, 1, 96, 96, 1, 96, 96, 1, 
    1, 96, 1, 96, 1, 96, 96, 1, 92, 1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 94, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 288, 1, 1, 96, 1, 96, 1, 
    95, 96, 1, 1, 96, 1, 96, 96, 1, 96, 288, 1, 288, 1, 288, 1, 288, 1, 288, 
    1, 96, 1, 1, 96, 288, 1, 1, 1, 288, 1, 1, 1, 1, 96, 1, 1, 288, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 288, 1, 288, 1, 288, 1, 1, 1, 1, 288, 1, 1, 1, 
    96, 288, 1, 1, 1, 1, 96, 1, 1, 288, 1, 288, 1, 96, 288, 1, 1, 1, 1, 96, 
    265, 1, 1, 1, 96, 288, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 288, 1, 1, 288, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 
    96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 96, 1, 1, 
    1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 288, 1, 1, 1, 1, 
    96, 288, 1, 1, 95, 1, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 288, 1, 1, 96, 1, 1, 
    1, 288, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 96, 1, 1, 95, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 66, 
    1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 96, 288, 1, 288, 1, 288, 1, 96, 1, 288, 1, 288, 
    288, 1, 288, 1, 96, 1, 288, 1, 288, 1, 288, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 48, 48, 1, 96, 1, 
    1, 1, 24, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 288, 1, 
    288, 1, 288, 1, 288, 1, 96, 1, 1, 288, 288, 1, 288, 1, 288, 1, 288, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 288, 
    288, 1, 288, 1, 1, 288, 288, 1, 288, 288, 1, 288, 1, 288, 288, 1, 288, 
    288, 1, 288, 288, 1, 288, 288, 288, 1, 288, 1, 288, 1, 1, 288, 1, 288, 
    288, 1, 288, 1, 288, 1, 288, 1, 1, 288, 288, 288, 288, 1, 288, 1, 288, 
    288, 1, 288, 1, 96, 1, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 
    1, 1, 1, 24, 96, 1, 96, 1, 96, 1, 1, 1, 1, 24, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 24, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 96, 96, 96, 96, 96, 1, 96, 96, 24, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 96, 96, 93, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 96, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    96, 96, 1, 1, 96, 96, 96, 1, 1, 96, 1, 1, 1, 96, 24, 1, 96, 1, 96, 1, 96, 
    1, 1, 24, 1, 24, 1, 1, 96, 24, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 95, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 91, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 24, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 72, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 95, 1, 1, 96, 1, 1, 95, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 94, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 94, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 73, 
    1, 1, 1, 96, 96, 1, 24, 1, 1, 96, 1, 96, 48, 1, 1, 24, 1, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 95, 1, 1, 94, 96, 1, 1, 96, 
    1, 96, 84, 1, 1, 1, 1, 96, 1, 48, 1, 48, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 48, 1, 24, 1, 24, 1, 24, 24, 1, 96, 96, 24, 24, 24, 24, 96, 96, 
    1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 24, 1, 24, 24, 48, 48, 1, 1, 96, 24, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 24, 1, 24, 96, 1, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 24, 1, 48, 96, 96, 1, 1, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 24, 24, 1, 96, 96, 1, 
    96, 1, 48, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 24, 1, 
    1, 48, 1, 1, 24, 24, 1, 24, 48, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 221, 92, 1, 96, 1, 89, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 24, 24, 96, 96, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    264, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 95, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 95, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 96, 
    1, 95, 94, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 96, 96, 96, 1, 
    96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 203, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 24, 1, 24, 1, 24, 1, 92, 1, 24, 1, 24, 95, 1, 1, 96, 96, 1, 1, 96, 1, 
    96, 24, 1, 1, 48, 1, 48, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 96, 1, 96, 96, 96, 1, 96, 96, 1, 96, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 1, 24, 1, 24, 24, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 24, 96, 1, 1, 96, 1, 92, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 24, 96, 1, 96, 1, 1, 1, 96, 1, 1, 24, 24, 1, 1, 24, 96, 
    1, 1, 1, 24, 1, 96, 1, 24, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 96, 1, 1, 1, 1, 1, 
    1, 24, 1, 24, 24, 1, 24, 1, 23, 1, 24, 24, 1, 96, 1, 24, 96, 96, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 24, 96, 1, 1, 1, 96, 1, 1, 24, 1, 1, 96, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 24, 24, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 91, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 95, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 95, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 92, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 93, 1, 1, 96, 1, 96, 1, 1, 1, 1, 92, 1, 96, 1, 1, 
    24, 1, 96, 1, 96, 1, 24, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 94, 1, 1, 92, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 48, 1, 1, 24, 1, 1, 
    96, 48, 1, 1, 48, 1, 24, 1, 1, 1, 96, 1, 1, 23, 1, 48, 1, 24, 24, 1, 96, 
    1, 1, 1, 24, 48, 1, 1, 24, 48, 1, 1, 48, 1, 96, 96, 1, 96, 1, 1, 48, 1, 
    48, 1, 96, 1, 48, 1, 96, 96, 1, 1, 1, 48, 1, 48, 1, 96, 1, 24, 1, 48, 96, 
    1, 96, 1, 1, 96, 96, 1, 1, 96, 48, 1, 1, 48, 1, 48, 1, 1, 96, 1, 96, 1, 
    48, 1, 48, 1, 96, 1, 24, 1, 96, 48, 1, 48, 96, 1, 48, 1, 1, 48, 1, 1, 96, 
    1, 1, 56, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 
    95, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 95, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 48, 1, 48, 48, 1, 
    48, 48, 48, 96, 1, 1, 48, 1, 48, 48, 1, 48, 1, 48, 1, 48, 1, 1, 48, 96, 
    1, 1, 96, 96, 1, 1, 48, 48, 1, 48, 48, 48, 1, 1, 48, 1, 95, 1, 96, 1, 1, 
    1, 48, 1, 48, 1, 48, 1, 47, 96, 1, 96, 1, 1, 24, 48, 48, 1, 1, 1, 24, 1, 
    48, 96, 1, 48, 24, 1, 24, 1, 48, 24, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 
    1, 24, 24, 1, 48, 24, 1, 24, 1, 24, 96, 1, 1, 24, 24, 96, 1, 96, 1, 96, 
    1, 24, 1, 1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 24, 24, 1, 96, 96, 1, 96, 
    24, 24, 96, 1, 1, 24, 24, 1, 24, 1, 96, 96, 96, 1, 1, 24, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 1, 48, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 288, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 96, 
    1, 1, 96, 96, 1, 24, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 96, 1, 90, 94, 1, 
    48, 96, 1, 23, 24, 1, 48, 24, 48, 1, 96, 1, 24, 1, 48, 1, 48, 1, 93, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 25, 1, 96, 1, 93, 1, 1, 1, 
    95, 1, 96, 1, 82, 1, 96, 1, 96, 81, 1, 96, 96, 1, 96, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 24, 48, 1, 48, 1, 48, 1, 96, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 91, 1, 1, 96, 96, 96, 96, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 95, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 96, 96, 96, 96, 1, 1, 96, 2, 96, 1, 1, 96, 96, 96, 1, 96, 1, 1, 96, 
    1, 96, 89, 1, 1, 1, 48, 1, 1, 1, 96, 96, 1, 96, 96, 1, 1, 48, 1, 1, 48, 
    1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 76, 36, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 24, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 48, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 96, 96, 1, 96, 1, 1, 1, 48, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 93, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 
    96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 95, 96, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 94, 95, 92, 96, 96, 1, 96, 96, 96, 1, 1, 96, 48, 48, 48, 96, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 48, 1, 1, 
    95, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 96, 48, 48, 1, 1, 96, 96, 96, 1, 
    95, 1, 1, 96, 1, 1, 1, 95, 48, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 48, 1, 84, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 96, 1, 1, 1, 96, 96, 
    96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 288, 1, 96, 1, 1, 96, 1, 
    1, 96, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 288, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 96, 94, 1, 96, 
    96, 96, 1, 1, 85, 88, 1, 96, 1, 96, 48, 1, 48, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 48, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 48, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 94, 
    1, 24, 96, 1, 42, 43, 1, 1, 96, 288, 1, 96, 1, 44, 40, 1, 96, 1, 1, 288, 
    1, 1, 96, 96, 1, 1, 96, 1, 96, 95, 1, 47, 48, 1, 96, 1, 1, 96, 48, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 48, 1, 48, 1, 96, 1, 48, 1, 48, 1, 
    48, 96, 1, 1, 48, 48, 1, 48, 48, 1, 95, 48, 89, 48, 48, 48, 48, 1, 96, 1, 
    48, 48, 48, 48, 48, 1, 48, 48, 1, 48, 1, 96, 48, 1, 48, 48, 96, 1, 48, 1, 
    48, 24, 1, 1, 48, 96, 1, 1, 96, 48, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 48, 1, 48, 48, 1, 96, 48, 1, 63, 1, 96, 1, 48, 1, 1, 96, 1, 96, 
    48, 48, 1, 48, 1, 48, 1, 48, 1, 96, 96, 1, 96, 1, 48, 1, 96, 1, 48, 48, 
    96, 1, 48, 1, 48, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 69, 1, 48, 1, 
    1, 48, 33, 1, 96, 96, 1, 1, 1, 96, 1, 48, 96, 1, 96, 1, 48, 1, 1, 96, 96, 
    1, 95, 96, 1, 1, 1, 96, 1, 48, 1, 1, 96, 1, 1, 96, 48, 1, 1, 48, 1, 96, 
    1, 48, 1, 93, 1, 48, 1, 96, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 96, 96, 1, 96, 96, 1, 48, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 96, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 48, 1, 20, 1, 96, 1, 96, 1, 96, 
    48, 1, 48, 1, 1, 48, 48, 1, 1, 48, 1, 48, 46, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 48, 48, 1, 47, 48, 48, 1, 1, 40, 48, 1, 1, 48, 
    48, 1, 96, 48, 42, 1, 1, 1, 48, 1, 1, 47, 1, 1, 1, 47, 1, 96, 48, 96, 1, 
    48, 1, 48, 1, 1, 48, 1, 1, 96, 1, 1, 1, 48, 1, 48, 1, 48, 1, 1, 48, 48, 
    1, 48, 1, 96, 1, 48, 1, 1, 96, 1, 48, 1, 1, 48, 48, 1, 48, 48, 48, 1, 47, 
    1, 48, 48, 1, 48, 1, 1, 46, 96, 1, 48, 1, 1, 24, 96, 1, 1, 96, 1, 48, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 48, 1, 48, 24, 1, 96, 1, 96, 
    1, 1, 96, 24, 1, 96, 1, 96, 1, 288, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 97, 96, 1, 96, 1, 48, 1, 96, 
    92, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 48, 1, 96, 1, 1, 96, 95, 96, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 288, 1, 
    1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 288, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 288, 1, 1, 288, 1, 1, 264, 1, 1, 96, 1, 95, 1, 1, 1, 92, 
    1, 96, 1, 1, 96, 1, 96, 96, 96, 1, 1, 1, 96, 1, 288, 1, 1, 288, 1, 1, 96, 
    1, 96, 1, 288, 1, 1, 288, 1, 1, 288, 1, 288, 1, 1, 1, 288, 1, 1, 1, 288, 
    1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    96, 144, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 288, 1, 1, 93, 1, 96, 1, 1, 1, 1, 92, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 96, 1, 1, 
    96, 96, 1, 1, 96, 288, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 288, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 96, 288, 1, 1, 96, 1, 96, 96, 96, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 95, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 96, 96, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 
    96, 24, 24, 24, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 92, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 
    24, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 24, 24, 1, 
    90, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 
    96, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 95, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 
    96, 1, 96, 1, 96, 96, 1, 96, 95, 1, 1, 96, 96, 1, 95, 95, 48, 1, 1, 48, 
    1, 1, 48, 1, 1, 1, 96, 1, 1, 48, 1, 48, 1, 1, 48, 48, 1, 1, 48, 1, 48, 1, 
    48, 1, 48, 1, 1, 1, 92, 1, 96, 1, 1, 1, 48, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    48, 48, 1, 1, 1, 48, 1, 1, 91, 1, 48, 48, 1, 1, 48, 1, 1, 1, 48, 1, 48, 
    1, 1, 48, 1, 288, 1, 97, 1, 95, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 96, 1, 
    96, 96, 287, 1, 1, 48, 1, 96, 1, 97, 1, 1, 1, 1, 1, 96, 288, 1, 1, 288, 
    94, 1, 1, 1, 96, 288, 1, 97, 1, 96, 1, 1, 97, 96, 1, 96, 1, 48, 1, 96, 
    96, 1, 1, 96, 1, 1, 1, 48, 1, 43, 1, 1, 48, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 48, 1, 48, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 
    1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 48, 96, 1, 1, 96, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 48, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 48, 96, 48, 1, 
    288, 1, 288, 1, 96, 288, 1, 288, 1, 1, 288, 1, 93, 288, 1, 288, 1, 288, 
    1, 288, 1, 1, 288, 1, 288, 288, 1, 1, 288, 1, 288, 1, 96, 1, 96, 96, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 48, 1, 96, 1, 90, 
    96, 96, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 48, 1, 48, 1, 95, 96, 1, 96, 
    1, 1, 96, 1, 48, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 48, 1, 48, 1, 96, 96, 1, 48, 1, 1, 1, 96, 1, 1, 96, 1, 1, 95, 
    288, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 93, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 95, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 24, 96, 1, 1, 96, 1, 1, 22, 1, 96, 1, 24, 24, 1, 
    96, 1, 96, 1, 96, 96, 1, 24, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 94, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 49, 96, 1, 1, 1, 1, 96, 
    288, 48, 1, 1, 288, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    9, 96, 1, 288, 1, 288, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 24, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 288, 1, 96, 288, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 288, 1, 1, 1, 1, 96, 1, 1, 1, 288, 
    96, 1, 135, 1, 1, 1, 96, 1, 288, 1, 141, 96, 1, 1, 34, 1, 1, 1, 1, 95, 1, 
    1, 96, 288, 1, 1, 96, 1, 96, 1, 1, 1, 93, 1, 1, 1, 96, 288, 1, 288, 1, 1, 
    1, 288, 1, 1, 96, 1, 1, 288, 1, 1, 1, 1, 288, 1, 1, 288, 1, 1, 1, 24, 1, 
    1, 24, 1, 1, 1, 96, 288, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 288, 264, 1, 1, 287, 1, 1, 1, 1, 96, 96, 96, 1, 96, 1, 96, 
    288, 1, 96, 96, 1, 96, 273, 1, 96, 1, 96, 1, 1, 96, 24, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 24, 24, 96, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 48, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 92, 1, 96, 1, 96, 96, 
    96, 1, 96, 1, 96, 96, 1, 1, 120, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 105, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 
    1, 1, 92, 1, 96, 1, 1, 96, 240, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 96, 1, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 120, 240, 96, 1, 120, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 
    45, 1, 1, 1, 1, 240, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 288, 1, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 
    1, 48, 1, 24, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 95, 1, 48, 
    48, 1, 1, 1, 97, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 96, 1, 96, 1, 48, 1, 1, 96, 96, 1, 93, 1, 1, 1, 1, 48, 1, 
    48, 48, 1, 48, 1, 1, 48, 1, 96, 48, 1, 96, 1, 1, 96, 1, 48, 1, 96, 1, 96, 
    1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 48, 1, 96, 288, 1, 1, 96, 1, 48, 1, 96, 
    1, 96, 1, 96, 1, 288, 1, 96, 1, 96, 1, 288, 1, 1, 96, 1, 1, 48, 1, 288, 
    96, 1, 288, 144, 1, 96, 1, 1, 1, 48, 1, 48, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 99, 1, 99, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 48, 1, 96, 1, 97, 96, 1, 1, 96, 1, 96, 48, 1, 
    96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 94, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 98, 96, 96, 1, 
    96, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 288, 1, 288, 1, 1, 96, 1, 94, 1, 96, 96, 1, 96, 96, 1, 96, 1, 
    81, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 
    96, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 
    1, 96, 96, 96, 96, 1, 96, 96, 96, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 
    1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 96, 1, 96, 1, 26, 1, 96, 96, 96, 1, 
    96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 96, 96, 1, 
    96, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 96, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 18, 1, 96, 1, 96, 1, 95, 1, 1, 1, 96, 96, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 96, 96, 1, 96, 96, 96, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 
    96, 96, 96, 1, 96, 1, 89, 96, 1, 96, 96, 1, 1, 96, 92, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 
    1, 96, 48, 1, 48, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 96, 1, 96, 96, 96, 1, 96, 96, 1, 24, 96, 1, 96, 96, 1, 1, 
    96, 96, 1, 96, 1, 96, 1, 96, 1, 48, 1, 1, 96, 1, 48, 1, 96, 96, 1, 96, 1, 
    96, 1, 25, 1, 25, 96, 96, 1, 88, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 96, 1, 1, 47, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 96, 1, 1, 96, 96, 96, 1, 1, 96, 96, 96, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 82, 1, 96, 1, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 96, 96, 
    96, 1, 1, 1, 96, 92, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 14, 96, 1, 1, 1, 24, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 95, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 
    96, 96, 96, 96, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    288, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 88, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 
    1, 87, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 96, 96, 1, 144, 96, 1, 1, 144, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 288, 1, 96, 1, 96, 1, 1, 96, 1, 288, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 288, 96, 288, 1, 1, 96, 1, 1, 288, 1, 1, 96, 1, 1, 1, 288, 1, 
    1, 96, 1, 1, 1, 189, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 144, 1, 96, 1, 96, 1, 96, 1, 288, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 
    1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 90, 1, 96, 1, 96, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 95, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 96, 96, 1, 96, 1, 96, 1, 96, 1, 81, 1, 96, 1, 
    96, 1, 96, 96, 1, 82, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 96, 88, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 86, 96, 1, 1, 96, 37, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 94, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 90, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 92, 1, 96, 96, 
    1, 1, 1, 96, 8, 1, 1, 96, 1, 96, 1, 96, 1, 144, 1, 96, 1, 58, 96, 1, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 48, 1, 96, 48, 
    1, 1, 1, 48, 96, 1, 47, 1, 1, 1, 46, 48, 1, 1, 48, 1, 48, 1, 48, 1, 48, 
    1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 96, 1, 48, 1, 288, 1, 1, 288, 1, 1, 96, 
    1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 95, 1, 95, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 95, 96, 288, 1, 1, 96, 
    96, 1, 96, 288, 1, 1, 96, 1, 288, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 288, 288, 288, 288, 
    288, 96, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1440, 1, 1, 1, 
    288, 96, 96, 1, 48, 1, 96, 96, 1, 1, 288, 1, 1, 1, 278, 96, 1, 96, 1, 1, 
    288, 1, 288, 1, 288, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 96, 96, 1, 96, 1, 288, 1, 96, 1, 1, 96, 96, 51, 95, 
    1, 1, 96, 1, 1, 96, 1, 96, 96, 96, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    24, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 96, 1, 1, 
    96, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 288, 1, 288, 1, 96, 1, 75, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 24, 24, 1, 190, 1, 1, 
    96, 1, 47, 48, 1, 48, 1, 96, 1, 286, 96, 1, 1, 96, 1, 1, 96, 93, 1, 96, 
    1, 96, 1, 94, 1, 1, 48, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 96, 1, 96, 95, 1, 96, 1, 96, 1, 1, 95, 1, 96, 1, 96, 1, 96, 
    46, 96, 1, 96, 48, 1, 96, 48, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 
    1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 93, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 69, 1, 49, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 
    76, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 95, 
    1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 62, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 34, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 35, 
    1, 1, 86, 1, 96, 96, 1, 1, 96, 1, 96, 1, 95, 1, 96, 88, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 94, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 50, 
    96, 1, 1, 96, 1, 96, 1, 73, 96, 1, 1, 57, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 95, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 
    37, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 95, 
    96, 1, 95, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 93, 1, 96, 1, 96, 1, 
    92, 1, 84, 1, 32, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 96, 1, 
    96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 288, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 288, 1, 1, 288, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 88, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 288, 1, 1, 
    1, 288, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 95, 1, 96, 
    1, 1, 96, 1, 1, 96, 96, 96, 94, 88, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 96, 96, 1, 96, 62, 62, 1, 96, 1, 1, 89, 1, 96, 1, 1, 96, 1, 1, 
    92, 1, 96, 1, 96, 96, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    87, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 95, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 14, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 289, 1, 96, 288, 96, 96, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 25, 1, 1, 96, 96, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 1, 84, 1, 
    96, 1, 96, 1, 38, 1, 91, 1, 99, 1, 96, 1, 81, 1, 95, 1, 33, 1, 1, 97, 1, 
    1, 94, 1, 91, 1, 93, 1, 1, 94, 1, 89, 1, 1, 88, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 88, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 288, 288, 1, 288, 
    1, 1, 96, 1, 1, 1, 288, 1, 288, 288, 1, 288, 1, 288, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 96, 1, 288, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 
    288, 1, 288, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 145, 1, 288, 267, 1, 96, 
    1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 1, 1, 29, 94, 1, 1, 96, 89, 1, 1, 96, 96, 1, 1, 95, 1, 96, 1, 96, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 95, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 96, 96, 1, 1, 96, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 90, 1, 96, 1, 71, 
    1, 1, 95, 1, 1, 96, 96, 96, 1, 96, 1, 96, 1, 52, 1, 1, 96, 96, 1, 96, 96, 
    1, 1, 96, 49, 1, 95, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 288, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 288, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    96, 96, 1, 96, 96, 1, 96, 80, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 94, 96, 1, 96, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 94, 96, 1, 1, 96, 1, 1, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 96, 1, 95, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 92, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 
    1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 96, 45, 96, 1, 1, 96, 81, 
    1, 96, 1, 1, 96, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 24, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 88, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 90, 288, 1, 288, 4, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 94, 1, 83, 96, 96, 1, 96, 1, 1, 1, 96, 89, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 92, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 69, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 54, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 36, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 1, 94, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 97, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 1, 94, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 288, 1, 288, 1, 1, 288, 1, 264, 1, 1, 
    1, 92, 288, 1, 1, 1, 96, 288, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 288, 288, 1, 288, 1, 1, 288, 1, 288, 1, 1, 1, 288, 1, 24, 
    1, 1, 1, 281, 1, 288, 1, 1, 288, 1, 287, 1, 288, 1, 288, 1, 288, 1, 1, 
    24, 1, 1, 288, 285, 1, 288, 1, 288, 264, 1, 288, 1, 288, 1, 288, 1, 1, 
    288, 288, 1, 288, 264, 1, 290, 1, 1, 288, 288, 1, 1, 288, 1, 1, 96, 48, 
    1, 1, 96, 1, 1, 1, 48, 1, 1, 96, 47, 1, 1, 48, 1, 96, 48, 1, 1, 1, 94, 
    48, 1, 1, 1, 264, 288, 1, 48, 1, 288, 1, 288, 1, 1, 288, 1, 288, 1, 1, 
    255, 287, 1, 48, 1, 96, 1, 46, 1, 1, 1, 1, 96, 96, 46, 1, 1, 1, 96, 94, 
    1, 1, 96, 1, 24, 24, 1, 96, 1, 96, 1, 46, 24, 1, 96, 96, 1, 96, 1, 96, 
    48, 1, 24, 24, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    1, 48, 24, 1, 96, 1, 61, 1, 96, 1, 48, 48, 1, 48, 1, 48, 1, 24, 1, 48, 1, 
    1, 1, 24, 1, 1, 96, 277, 1, 1, 1, 1, 89, 1, 24, 288, 1, 1, 288, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 288, 1, 96, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 22, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 98, 96, 1, 1, 47, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 92, 1, 1, 1, 1, 55, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 24, 96, 1, 1, 24, 24, 1, 
    286, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 
    156, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 96, 1, 96, 1, 1, 1, 85, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 86, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 96, 96, 96, 96, 1, 96, 1, 96, 96, 96, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 96, 1, 24, 1, 1, 1, 24, 1, 1, 
    1, 24, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 
    1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 1, 48, 48, 1, 
    1, 96, 1, 48, 1, 1, 24, 1, 1, 1, 48, 96, 1, 1, 1, 48, 1, 96, 1, 96, 48, 
    1, 1, 48, 1, 1, 48, 1, 24, 1, 24, 1, 96, 1, 1, 1, 48, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 24, 1, 1, 48, 1, 1, 96, 1, 92, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 24, 24, 96, 1, 96, 1, 1, 96, 48, 1, 1, 96, 1, 
    48, 1, 1, 48, 1, 96, 1, 1, 48, 1, 1, 96, 1, 1, 26, 1, 1, 1, 1, 96, 1, 96, 
    1, 48, 1, 48, 1, 1, 1, 96, 84, 48, 1, 1, 24, 95, 1, 24, 1, 96, 96, 1, 1, 
    96, 96, 96, 1, 70, 1, 48, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    24, 1, 1, 96, 1, 24, 1, 1, 96, 1, 1, 48, 24, 1, 1, 96, 96, 1, 1, 92, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 94, 1, 96, 1, 1, 24, 1, 1, 96, 1, 
    1, 48, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 23, 
    1, 96, 1, 48, 1, 1, 96, 1, 1, 94, 1, 1, 48, 1, 1, 96, 1, 1, 1, 1, 48, 1, 
    48, 1, 1, 96, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 96, 1, 96, 1, 96, 288, 
    1, 1, 96, 1, 1, 1, 1, 290, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 24, 1, 
    1, 1, 96, 96, 1, 1, 96, 1, 48, 1, 1, 96, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 
    48, 1, 96, 1, 1, 1, 48, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 92, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 288, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 48, 48, 1, 1, 48, 48, 1, 1, 24, 
    1, 288, 24, 1, 48, 1, 48, 1, 96, 1, 1, 1, 48, 1, 48, 1, 1, 96, 1, 1, 1, 
    48, 1, 1, 96, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 24, 1, 24, 1, 48, 1, 1, 
    48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 96, 24, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 48, 1, 1, 48, 1, 24, 1, 1, 48, 1, 1, 1, 48, 48, 1, 96, 
    1, 1, 48, 1, 1, 96, 96, 1, 48, 1, 48, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 24, 24, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 93, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 24, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    73, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 24, 24, 1, 24, 96, 1, 1, 1, 288, 1, 96, 1, 1, 96, 1, 96, 
    96, 24, 30, 1, 24, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 92, 1, 
    96, 96, 1, 24, 1, 96, 24, 1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 24, 27, 90, 15, 1, 1, 96, 1, 24, 24, 1, 1, 96, 24, 1, 96, 1, 96, 
    1, 96, 1, 24, 96, 1, 1, 1, 1, 96, 1, 1, 86, 1, 1, 60, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 62, 1, 96, 1, 1, 96, 1, 1, 96, 1, 48, 1, 1, 
    1, 48, 48, 1, 1, 24, 1, 1, 96, 1, 48, 1, 1, 48, 1, 1, 1, 48, 1, 48, 1, 1, 
    1, 96, 96, 1, 1, 1, 48, 1, 96, 1, 1, 48, 1, 48, 1, 1, 48, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 62, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 93, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 48, 
    1, 1, 1, 1, 37, 48, 1, 1, 96, 1, 1, 24, 1, 1, 96, 1, 1, 48, 1, 1, 1, 48, 
    1, 48, 1, 1, 96, 1, 1, 95, 1, 1, 96, 1, 1, 24, 1, 96, 1, 48, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 48, 96, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 24, 144, 1, 
    1, 1, 24, 1, 23, 96, 1, 1, 1, 24, 48, 1, 1, 48, 96, 1, 1, 48, 1, 24, 1, 
    96, 1, 1, 46, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 48, 1, 48, 1, 24, 1, 48, 
    1, 1, 24, 1, 1, 1, 1, 48, 96, 24, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 24, 1, 
    24, 1, 1, 48, 1, 1, 1, 1, 24, 1, 96, 1, 1, 96, 88, 48, 1, 1, 48, 1, 1, 
    48, 1, 1, 48, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 90, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 48, 1, 96, 96, 96, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 24, 48, 96, 96, 
    23, 24, 24, 1, 96, 1, 46, 48, 96, 96, 48, 24, 24, 24, 96, 1, 48, 96, 48, 
    288, 96, 96, 1, 96, 24, 1, 48, 48, 1, 48, 48, 48, 24, 1, 96, 96, 96, 1, 
    1, 1, 1, 96, 1, 1, 285, 288, 1, 1, 288, 1, 1, 96, 1, 96, 96, 1, 1, 288, 
    1, 1, 96, 1, 1, 1, 288, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 24, 1, 
    1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 95, 1, 96, 1, 
    1, 1, 96, 1, 24, 24, 1, 96, 1, 1, 1, 50, 1, 1, 1, 96, 1, 1, 48, 96, 1, 1, 
    1, 48, 48, 48, 24, 24, 1, 1, 24, 96, 1, 48, 48, 1, 96, 1, 48, 1, 1, 48, 
    48, 1, 48, 48, 1, 48, 24, 96, 1, 1, 1, 1, 96, 48, 48, 48, 1, 96, 1, 96, 
    1, 96, 96, 1, 1, 1, 24, 24, 96, 1, 1, 1, 48, 1, 1, 24, 1, 1, 48, 24, 1, 
    1, 240, 1, 1, 1, 1, 24, 1, 1, 96, 24, 96, 1, 96, 56, 1, 96, 1, 48, 1, 96, 
    1, 96, 1, 96, 1, 48, 1, 1, 1, 1, 96, 48, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 48, 1, 96, 1, 1, 96, 1, 48, 1, 1, 48, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 48, 1, 96, 1, 48, 1, 1, 48, 96, 48, 1, 48, 1, 1, 1, 1, 96, 1, 
    96, 1, 96, 96, 1, 96, 4, 1, 96, 96, 1, 96, 1, 96, 1, 96, 48, 1, 48, 1, 
    48, 96, 1, 1, 48, 1, 1, 96, 48, 1, 48, 1, 1, 1, 33, 1, 48, 48, 1, 48, 1, 
    48, 1, 48, 1, 96, 1, 96, 96, 1, 36, 1, 1, 1, 24, 1, 1, 24, 1, 1, 240, 1, 
    1, 1, 1, 96, 24, 1, 1, 24, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 96, 96, 96, 1, 
    1, 1, 1, 1, 240, 1, 1, 24, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 96, 1, 
    1, 1, 96, 1, 1, 56, 1, 24, 96, 48, 48, 1, 1, 96, 96, 48, 1, 96, 1, 96, 
    96, 240, 96, 1, 1, 48, 96, 1, 48, 48, 96, 1, 96, 96, 1, 96, 48, 1, 48, 
    96, 1, 1, 1, 1, 48, 1, 96, 240, 1, 1, 1, 1, 24, 1, 1, 1, 48, 1, 48, 1, 1, 
    1, 40, 1, 1, 48, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 96, 1, 48, 1, 1, 1, 
    24, 1, 1, 1, 1, 24, 1, 1, 24, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 95, 1, 1, 96, 96, 1, 85, 1, 1, 1, 96, 1, 48, 1, 96, 1, 
    1, 1, 1, 90, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 95, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 73, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 72, 1, 96, 
    96, 1, 94, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 94, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 95, 1, 96, 1, 
    96, 96, 1, 96, 96, 1, 1, 1, 1, 95, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 87, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 
    96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 60, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 90, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 95, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 95, 
    1, 1, 288, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 288, 1, 1, 1, 1, 95, 96, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 288, 1, 1, 1, 96, 1, 1, 1, 96, 1, 288, 288, 288, 
    1, 288, 288, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    95, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 288, 1, 1, 288, 1, 1, 95, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    288, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 
    1, 96, 1, 96, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 
    1, 95, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 288, 1, 288, 1, 1, 1, 96, 1, 1, 
    288, 1, 1, 288, 1, 1, 96, 1, 96, 1, 288, 1, 1, 288, 1, 1, 96, 1, 288, 1, 
    288, 1, 288, 1, 288, 1, 288, 1, 288, 1, 288, 1, 288, 288, 1, 1, 96, 1, 1, 
    288, 1, 288, 1, 1, 288, 288, 1, 288, 1, 1, 288, 288, 1, 288, 1, 288, 1, 
    1, 1, 1, 1, 288, 1, 288, 1, 288, 1, 288, 1, 1, 196, 288, 1, 1, 288, 288, 
    1, 1, 288, 288, 1, 1, 288, 1, 288, 1, 288, 1, 288, 1, 288, 288, 1, 288, 
    96, 1, 1, 288, 1, 288, 1, 1, 288, 288, 1, 1, 96, 96, 1, 1, 96, 96, 96, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 93, 1, 96, 1, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 95, 1, 
    96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 68, 1, 1, 96, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    96, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 92, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 95, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 46, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 11, 96, 1, 
    1, 288, 1, 96, 1, 1, 96, 1, 1, 96, 1, 288, 1, 288, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 93, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 16, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 96, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 144, 1, 1, 1, 
    96, 1, 288, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 95, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 
    1, 1, 64, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 288, 288, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 80, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 93, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 93, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 288, 96, 1, 1, 96, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 94, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 94, 1, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 96, 1, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 90, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 91, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 96, 1, 96, 1, 94, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    101, 1, 101, 1, 93, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 94, 
    96, 1, 1, 1, 96, 1, 96, 1, 23, 1, 1, 96, 94, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 95, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 95, 1, 96, 96, 96, 
    1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 192, 96, 1, 192, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 94, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 95, 96, 1, 96, 1, 96, 1, 96, 96, 96, 96, 1, 
    96, 1, 96, 1, 81, 1, 96, 1, 44, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 65, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 119, 1, 
    1, 96, 1, 95, 1, 1, 96, 1, 96, 1, 48, 98, 98, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 95, 1, 164, 1, 164, 1, 96, 1, 
    96, 1, 1, 94, 97, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 100, 1, 96, 1, 1, 96, 1, 99, 
    1, 96, 96, 1, 1, 96, 1, 1, 97, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 97, 1, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 24, 24, 1, 
    24, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 94, 83, 1, 96, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 62, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    94, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 92, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 92, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 
    96, 1, 1, 96, 1, 96, 96, 1, 35, 1, 1, 43, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    96, 1, 96, 76, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    80, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 24, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 95, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    89, 1, 96, 1, 76, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 85, 1, 96, 1, 96, 
    1, 96, 1, 62, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 90, 96, 1, 96, 94, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    1, 96, 1, 95, 1, 96, 91, 1, 95, 96, 96, 1, 96, 1, 96, 1, 100, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 98, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 94, 1, 96, 
    1, 288, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 288, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 93, 1, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 49, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 94, 1, 1, 95, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 85, 1, 85, 1, 85, 1, 85, 85, 1, 1, 86, 1, 1, 82, 1, 82, 82, 1, 
    1, 1, 1, 82, 1, 82, 1, 82, 1, 86, 1, 1, 1, 96, 1, 96, 96, 1, 1, 86, 1, 
    86, 1, 86, 1, 1, 87, 1, 59, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 93, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 84, 1, 1, 1, 84, 1, 84, 1, 78, 96, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 35, 1, 40, 96, 1, 96, 1, 96, 1, 
    1, 1, 84, 1, 84, 1, 1, 84, 1, 1, 84, 1, 1, 1, 84, 1, 1, 1, 96, 1, 96, 96, 
    1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 84, 96, 1, 89, 1, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 1, 42, 1, 1, 96, 1, 96, 1, 96, 96, 96, 1, 96, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 96, 96, 1, 1, 96, 20, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 144, 1, 1, 1, 48, 1, 
    96, 1, 1, 96, 1, 1, 96, 227, 1, 1, 1, 48, 96, 96, 1, 1, 96, 1, 1, 1, 1, 
    144, 1, 144, 1, 144, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 91, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 53, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 96, 1, 48, 1, 96, 1, 96, 1, 1, 96, 1, 48, 1, 96, 96, 1, 96, 1, 
    96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 1, 96, 1, 96, 96, 
    1, 96, 1, 96, 96, 1, 96, 49, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 32, 1, 86, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 96, 96, 96, 48, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 24, 1, 96, 1, 24, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 24, 1, 48, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 96, 96, 1, 96, 96, 96, 1, 96, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 95, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    94, 1, 96, 1, 66, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 93, 1, 96, 96, 1, 96, 1, 96, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 56, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 288, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 97, 1, 96, 1, 1, 95, 1, 96, 96, 1, 96, 96, 97, 97, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 72, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 81, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 89, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 97, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 56, 84, 1, 1, 96, 1, 96, 96, 1, 
    1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 99, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 41, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 52, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 28, 28, 1, 96, 1, 96, 1, 1, 96, 1, 44, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 1, 86, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 48, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 
    1, 96, 1, 96, 96, 96, 1, 89, 1, 48, 1, 1, 1, 1, 48, 96, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 112, 1, 1, 96, 96, 1, 1, 1, 96, 1, 108, 1, 104, 1, 1, 98, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 67, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 97, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 114, 1, 
    1, 108, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 106, 1, 96, 1, 1, 1, 96, 
    1, 1, 112, 1, 96, 1, 1, 107, 1, 131, 1, 101, 1, 127, 1, 137, 1, 1, 126, 
    1, 128, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 94, 1, 1, 1, 96, 1, 96, 1, 1, 97, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 
    96, 1, 96, 1, 1, 288, 97, 1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    95, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    1, 96, 1, 96, 96, 96, 96, 1, 1, 48, 1, 96, 1, 1, 42, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 87, 1, 96, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 96, 96, 1, 1, 1, 88, 
    1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 51, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 24, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 64, 
    1, 64, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 96, 1, 96, 96, 1, 96, 
    1, 96, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 1, 94, 1, 96, 1, 96, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 113, 1, 96, 96, 1, 96, 1, 96, 96, 1, 225, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 112, 1, 96, 1, 102, 1, 100, 1, 96, 1, 96, 1, 288, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 52, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 96, 96, 96, 1, 1, 96, 91, 1, 1, 96, 1, 1, 1, 96, 96, 96, 96, 
    96, 96, 1, 1, 24, 24, 96, 96, 96, 96, 96, 96, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 96, 96, 96, 96, 96, 
    96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 1, 96, 1, 96, 96, 
    1, 96, 1, 96, 96, 96, 96, 96, 96, 96, 95, 96, 96, 96, 96, 96, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 
    1, 1, 24, 1, 1, 48, 48, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 48, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 48, 1, 48, 
    1, 24, 1, 1, 35, 1, 1, 186, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 24, 1, 96, 1, 1, 1, 1, 96, 48, 1, 1, 96, 96, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    91, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 84, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 58, 1, 48, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 137, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 88, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 71, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 288, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 96, 
    96, 1, 96, 1, 1, 1, 24, 24, 1, 1440, 1, 24, 24, 1, 24, 24, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 890, 1, 1, 96, 1, 1, 96, 
    1, 89, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 288, 1, 1211, 
    1, 1, 96, 1, 1, 1, 1, 96, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 88, 1, 96, 1, 96, 
    1, 1, 1, 1, 288, 288, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    95, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1 ;

 v00010_value =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 144, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 87, 1, 1, 1, 
    97, 1, 95, 1, 1, 1, 1, 1, 144, 1, 1, 1, 111, 1, 1, 1, 144, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 26, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 144, 
    1, 1, 1, 1, 144, 1, 1, 144, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 
    1, 1, 96, 1, 1, 144, 1, 1, 1, 1, 144, 1, 1, 144, 1, 1, 1, 1, 1, 144, 1, 
    144, 1, 1, 1, 1, 144, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 93, 1, 1, 1, 1, 1, 93, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 240, 1, 226, 1, 1, 1, 1, 
    1, 240, 1, 240, 1, 1, 1, 240, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 120, 1, 
    240, 1, 1, 1, 240, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 52, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 24, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 24, 1, 1, 1, 1, 1, 20, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 1, 
    24, 1, 1, 1, 24, 1, 1, 120, 1, 1, 1, 1, 1, 24, 23, 1, 1, 120, 1, 1, 1, 1, 
    120, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 24, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 24, 1, 20, 1, 24, 1, 24, 1, 24, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 
    48, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 27, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 47, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 25, 1, 1, 1, 48, 1, 1, 1, 1, 
    48, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 46, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 231, 1, 1, 240, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 208, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 48, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 96, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 
    1, 288, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 92, 92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 103, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 24, 24, 1, 1, 1, 24, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 96, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 13, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    84, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 95, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 93, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 95, 1, 1, 1, 1, 61, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 93, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 73, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 84, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 93, 1, 1, 95, 1, 1, 61, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    91, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 96, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 89, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 95, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 94, 1, 95, 1, 1, 95, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 61, 1, 61, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 82, 1, 1, 1, 1, 1, 94, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 91, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 32, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 93, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 14, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 90, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 84, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 36, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 92, 1, 1, 1, 
    94, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 95, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 48, 1, 1, 1, 24, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 24, 1, 1, 1, 1, 96, 1, 1, 24, 1, 24, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 24, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 24, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 70, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 91, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 288, 1, 1, 
    1, 289, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 34, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 
    289, 1, 1, 1, 1, 1, 1, 192, 1, 1, 1, 288, 1, 1, 1, 288, 1, 1, 1, 288, 1, 
    1, 24, 1, 1, 1, 24, 1, 1, 1, 288, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 24, 1, 1, 24, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    24, 1, 1, 24, 1, 1, 24, 24, 24, 24, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 276, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 120, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 289, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 46, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 76, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 3, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 78, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    86, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 288, 1, 1, 1, 1, 
    288, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 144, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 288, 1, 1, 1, 96, 1, 1, 1, 288, 1, 1, 96, 1, 1, 189, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 25, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 89, 1, 1, 1, 1, 1, 95, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1440, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    97, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 51, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 35, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 36, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 21, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 47, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    22, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 92, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    22, 1, 1, 11, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 276, 276, 276, 276, 276, 276, 276, 276, 1, 1, 
    276, 276, 276, 276, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 72, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 50, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 48, 1, 1, 23, 1, 1, 48, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 24, 1, 1, 25, 1, 1, 1, 
    1, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 24, 1, 1, 1, 1, 
    1, 24, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 48, 96, 1, 1, 96, 1, 1, 96, 1, 72, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    94, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 93, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 45, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 67, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 25, 1, 25, 1, 25, 1, 25, 1, 
    1, 1, 1, 1, 1, 1, 144, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 42, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 5, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 18, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 95, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 93, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 85, 1, 20, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 94, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 82, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 90, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 24, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 96, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 84, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    84, 1, 1, 1, 1, 1, 83, 1, 1, 1, 1, 1, 84, 1, 1, 1, 84, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 95, 1, 1, 1, 1, 144, 1, 1, 1, 1, 1, 1, 1, 96, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 24, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 78, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 73, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 
    1, 1, 1, 1, 1, 1, 98, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 86, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 97, 1, 1, 1, 1, 1, 1, 1, 1, 96, 114, 
    1, 1, 108, 1, 1, 1, 1, 96, 1, 1, 1, 1, 87, 1, 1, 106, 1, 1, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 113, 1, 107, 1, 1, 1, 1, 101, 1, 1, 1, 1, 1, 126, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 25, 
    1, 1, 1, 1, 1, 24, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 49, 1, 
    1, 1, 48, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 96, 1, 97, 1, 1, 96, 1, 1, 96, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 96, 1, 1, 1, 48, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 40, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 24, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 64, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 47, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    96, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 91, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 96, 96, 96, 96, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 25, 25, 25, 25, 25, 25, 25, 
    25, 25, 25, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 93, 1, 93, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 95, 1, 95, 1, 95, 24, 1, 24, 1, 1, 24, 1, 24, 1, 1, 1, 24, 
    1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 24, 1, 1, 24, 1, 1, 
    1, 48, 24, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 48, 1, 24, 1, 1, 96, 1, 24, 1, 
    24, 1, 24, 1, 24, 1, 1, 24, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 48, 1, 48, 1, 24, 1, 
    1, 60, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 48, 1, 48, 1, 96, 1, 1, 24, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 24, 1, 24, 94, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    49, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 96, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 18, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 
    48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 85, 85, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 88, 
    1, 1, 85, 1, 1, 23, 1, 19, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 24, 1, 
    24, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 92, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    720, 720, 720, 720, 720, 720, 720, 720, 720, 720, 720, 720, 720, 720, 
    720, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 24, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 24, 24, 1, 1, 24, 1, 1, 1, 24, 
    1, 1, 1, 24, 1, 24, 1, 24, 1, 95, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 96, 1, 1, 90, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 82, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 52, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 35, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 19, 1, 19, 19, 23, 21, 24, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    24, 1, 24, 1, 1, 24, 1, 24, 6, 1, 8, 1, 19, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 10, 10, 1, 1, 23, 1, 5, 1, 18, 18, 1, 19, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1 ;

 v00095_value =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 144, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 78, 1, 97, 1, 
    1, 1, 95, 1, 1, 1, 1, 1, 144, 1, 1, 1, 96, 1, 1, 1, 144, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    37, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 144, 1, 
    1, 1, 1, 144, 1, 1, 144, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 96, 
    1, 1, 1, 1, 144, 1, 1, 1, 1, 144, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 144, 
    1, 1, 144, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    93, 1, 1, 1, 1, 1, 93, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 240, 1, 226, 1, 1, 1, 1, 1, 240, 1, 
    240, 1, 1, 1, 240, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 120, 1, 240, 1, 1, 1, 
    240, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 24, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 27, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 46, 1, 1, 1, 1, 1, 47, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 25, 1, 1, 1, 48, 1, 1, 48, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 231, 1, 1, 240, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 205, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 288, 1, 1, 
    1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 92, 92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 48, 1, 1, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 84, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 95, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 92, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 58, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    93, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 73, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 84, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 
    1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 90, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 89, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 88, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 94, 1, 95, 1, 1, 1, 1, 95, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 60, 1, 61, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 86, 1, 1, 1, 1, 94, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 91, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 32, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    93, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 84, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 12, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 22, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 36, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 92, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 90, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 
    289, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 289, 1, 1, 
    1, 1, 1, 1, 192, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 288, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 276, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 120, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 289, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 46, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 84, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 
    1, 288, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 44, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 67, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 97, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 83, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 21, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 22, 1, 1, 11, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 88, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 44, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 
    1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    73, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 50, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 23, 1, 1, 48, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 24, 1, 1, 25, 1, 1, 1, 1, 1, 
    24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 24, 1, 1, 1, 24, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 
    1, 24, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    1, 1, 96, 48, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 93, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 44, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 69, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 25, 1, 25, 1, 25, 1, 25, 1, 1, 1, 
    1, 1, 1, 1, 144, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 5, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 18, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 85, 1, 13, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    82, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 90, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 84, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 84, 1, 1, 1, 1, 1, 83, 1, 1, 1, 1, 1, 84, 1, 1, 1, 84, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 41, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 25, 1, 1, 
    1, 1, 1, 24, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 49, 1, 1, 1, 
    48, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 50, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 52, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 96, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    91, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 93, 1, 92, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 95, 1, 95, 1, 95, 1, 1, 24, 1, 24, 24, 1, 1, 1, 24, 1, 1, 1, 
    24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 24, 1, 1, 24, 1, 
    1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 96, 1, 24, 
    1, 24, 1, 24, 1, 24, 1, 1, 24, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    60, 1, 1, 1, 1, 1, 24, 1, 1, 96, 48, 1, 48, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 24, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 96, 31, 1, 1, 1, 
    1, 24, 24, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 18, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    96, 1, 1, 85, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 88, 85, 1, 1, 23, 1, 19, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 24, 1, 24, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 92, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 24, 1, 1, 1, 24, 1, 24, 1, 24, 1, 95, 1, 24, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 88, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    82, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 24, 1, 24, 1, 1, 1, 1, 1, 6, 1, 8, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1 ;

 v00035_value =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 90, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 36, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 15, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 276, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 33, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 12, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 65, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 48, 48, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 56, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 48, 
    1, 1, 1, 1, 1, 1, 45, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 48, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 24, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 7, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 25, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    19, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 v00036_value =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 240, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 90, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 34, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 15, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 276, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 36, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    65, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 25, 25, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 52, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 44, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 24, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 716, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 24, 
    1, 24, 24, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 7, 1, 1, 1, 1, 1, 1, 1, 1, 1, 25, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 19, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 v00045_value =
  96, 45, 96, 96, 1, 96, 96, 24, 24, 96, 48, 48, 96, 96, 96, 96, 96, 96, 96, 
    96, 24, 96, 96, 96, 48, 96, 24, 144, 96, 48, 96, 96, 96, 96, 48, 24, 96, 
    96, 96, 96, 96, 96, 96, 96, 96, 96, 142, 96, 96, 96, 144, 96, 24, 96, 96, 
    96, 144, 96, 24, 96, 144, 96, 144, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 95, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 43, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    240, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 90, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 288, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 288, 
    1, 1, 1, 1, 96, 288, 1, 1, 96, 1, 1, 1, 288, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 95, 1, 1, 1, 1, 69, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 95, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 93, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 94, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 85, 1, 1, 1, 85, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 95, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 92, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 86, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 42, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 92, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 48, 1, 1, 48, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 96, 48, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 48, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 89, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 288, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 93, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 42, 1, 1, 
    96, 1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 24, 1, 96, 1, 1, 1, 288, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 1, 288, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 
    288, 1, 1, 264, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 288, 1, 1, 288, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 288, 
    1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 288, 1, 1, 93, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 
    1, 24, 1, 1, 1, 96, 1, 1, 24, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 288, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 92, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 48, 1, 1, 1, 48, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 
    48, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 
    1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 48, 1, 288, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 48, 1, 288, 1, 1, 1, 1, 1, 1, 1, 
    1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 48, 1, 1, 1, 43, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 48, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 288, 1, 1, 288, 1, 1, 288, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 288, 1, 288, 1, 1, 288, 1, 288, 288, 1, 96, 1, 1, 288, 1, 288, 1, 
    288, 1, 288, 288, 1, 288, 1, 1, 288, 288, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 288, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 135, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 7, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 
    95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 288, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 288, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 43, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 288, 1, 
    1, 288, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 95, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 68, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 89, 
    1, 1, 1, 77, 1, 91, 1, 96, 1, 1, 1, 89, 1, 92, 1, 1, 62, 1, 1, 95, 1, 93, 
    1, 93, 1, 1, 92, 1, 92, 1, 1, 93, 1, 1, 4, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 56, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 48, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 47, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 22, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 40, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 92, 1, 1, 1, 1, 54, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 279, 1, 1, 
    1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 288, 1, 1, 288, 1, 1, 1, 1, 1, 
    1, 288, 1, 1, 288, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 
    1, 1, 24, 1, 1, 1, 96, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 48, 1, 96, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 96, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 92, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 48, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 96, 1, 1, 96, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    96, 1, 1, 48, 1, 1, 48, 1, 1, 24, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 48, 1, 1, 96, 1, 1, 24, 1, 1, 96, 1, 48, 1, 1, 1, 48, 1, 48, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 
    1, 48, 1, 1, 1, 1, 96, 1, 96, 1, 1, 48, 1, 1, 96, 1, 1, 48, 1, 1, 48, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 24, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 88, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 24, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 92, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 44, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 48, 48, 1, 1, 1, 48, 1, 1, 24, 1, 
    1, 1, 1, 48, 1, 1, 48, 48, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 96, 1, 
    1, 1, 24, 24, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 96, 1, 24, 1, 1, 96, 1, 1, 
    96, 1, 24, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 24, 1, 1, 96, 1, 
    24, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 
    1, 1, 96, 1, 1, 24, 1, 1, 96, 1, 1, 48, 48, 1, 1, 1, 1, 48, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 24, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 1, 144, 1, 1, 23, 1, 1, 1, 1, 24, 1, 
    1, 1, 48, 1, 1, 1, 144, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 
    1, 96, 1, 1, 1, 48, 1, 1, 1, 1, 1, 24, 1, 1, 48, 1, 24, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 24, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 50, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 55, 1, 96, 1, 48, 1, 1, 1, 96, 1, 
    96, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 48, 1, 
    1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 48, 1, 96, 1, 96, 1, 96, 1, 96, 1, 48, 
    1, 96, 1, 1, 48, 1, 1, 1, 48, 1, 48, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 71, 1, 1, 96, 1, 96, 1, 96, 1, 1, 48, 1, 48, 1, 1, 1, 96, 1, 48, 96, 
    1, 1, 48, 1, 48, 1, 1, 1, 33, 1, 1, 48, 1, 48, 1, 48, 1, 48, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 56, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 88, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 95, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 95, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 95, 1, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 288, 1, 1, 288, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 1, 288, 1, 1, 1, 96, 1, 1, 288, 1, 1, 288, 1, 1, 96, 
    1, 1, 1, 288, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1378, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 
    288, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 29, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 31, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 92, 1, 
    1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 288, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 
    1, 80, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 94, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 118, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 98, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 92, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 44, 1, 1, 
    1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 
    1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    48, 1, 48, 1, 48, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 48, 
    1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 32, 1, 1, 48, 1, 1, 48, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 91, 288, 96, 96, 
    96, 96, 96, 96, 1, 96, 96, 1, 1, 96, 96, 96, 96, 96, 96, 1, 96, 96, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 
    96, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 274, 96, 96, 96, 
    1, 1, 96, 1, 1, 96, 96, 96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 
    96, 48, 1, 1, 96, 1, 1, 1, 96, 98, 288, 17, 288, 96, 96, 1, 96, 96, 96, 
    99, 96, 96, 96, 96, 96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 
    1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 96, 96, 1, 1, 24, 96, 96, 1, 96, 1, 96, 
    96, 126, 126, 1, 96, 126, 96, 96, 96, 72, 96, 96, 48, 96, 263, 1, 1, 1, 
    1, 1, 1, 264, 96, 96, 96, 96, 96, 96, 96, 288, 96, 288, 288, 288, 288, 
    288, 288, 288, 288, 288, 288, 288, 288, 288, 288, 288, 96, 96, 288, 288, 
    288, 288, 288, 288, 288, 288, 288, 288, 288, 288, 1, 1, 288, 288, 288, 
    288, 288, 48, 288, 288, 288, 288, 288, 288, 288, 288, 48, 288, 288, 288, 
    288, 288, 288, 288, 288, 288, 288, 288, 288, 288, 1, 1, 288, 288, 288, 
    288, 288, 288, 288, 288, 1, 1, 288, 288, 288, 288, 288, 288, 288, 96, 48, 
    288, 1, 96, 288, 288, 288, 96, 96, 1, 1, 288, 288, 288, 1, 1, 288, 288, 
    288, 1, 288, 288, 288, 288, 96, 288, 288, 288, 288, 288, 288, 288, 96, 1, 
    1, 1, 1, 96, 96, 1, 1, 288, 96, 1, 96, 96, 48, 288, 288, 1, 1, 1, 288, 1, 
    1, 96, 96, 96, 38, 96, 1, 96, 48, 96, 48, 1, 1, 96, 48, 48, 1, 48, 96, 1, 
    1, 48, 48, 48, 96, 48, 96, 48, 96, 48, 288, 96, 48, 96, 288, 48, 1, 1, 1, 
    288, 288, 1, 1, 1, 1, 1, 288, 1, 1, 48, 48, 96, 1, 1, 1, 1, 1, 1, 48, 1, 
    1, 1, 1, 1, 1, 1, 96, 48, 96, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 96, 
    96, 48, 1, 96, 1, 1, 48, 288, 1, 1, 1, 1, 288, 48, 1, 1, 1, 1, 48, 96, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 48, 48, 1, 1, 48, 288, 96, 
    96, 1, 1, 288, 1, 1, 1, 288, 288, 288, 149, 96, 96, 1, 1, 48, 96, 96, 96, 
    24, 288, 1, 1, 1, 1, 48, 24, 288, 96, 96, 48, 96, 96, 1, 1, 288, 48, 1, 
    1, 96, 48, 48, 96, 48, 96, 1, 1, 96, 96, 48, 1, 1, 1, 1, 96, 24, 96, 1, 
    1, 48, 1, 96, 1, 288, 288, 288, 288, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 24, 48, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 48, 96, 1, 24, 288, 1, 1, 96, 
    48, 1, 1, 288, 1, 1, 1, 1, 48, 96, 288, 288, 96, 1, 1, 288, 1, 1, 1, 1, 
    89, 96, 95, 1, 1, 1, 1, 1, 288, 1, 1, 96, 96, 96, 96, 1, 1, 48, 96, 96, 
    288, 1, 1, 24, 1, 1, 96, 1, 1, 1, 288, 1, 1, 48, 96, 96, 96, 48, 96, 96, 
    96, 96, 96, 1, 1, 96, 1, 1, 96, 96, 96, 96, 96, 96, 1, 96, 96, 96, 96, 
    96, 96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 
    96, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 96, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 96, 96, 96, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 2, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    96, 96, 1, 1, 1, 144, 96, 1, 1, 24, 288, 1, 1, 288, 1, 1, 48, 96, 1, 96, 
    96, 24, 48, 96, 96, 1, 96, 1, 1, 48, 1, 1, 1, 96, 96, 96, 48, 96, 96, 1, 
    1, 1, 1, 48, 1, 1, 48, 96, 55, 1, 1, 288, 288, 1, 288, 288, 96, 288, 149, 
    96, 1, 1, 48, 288, 288, 288, 288, 48, 48, 1, 1, 273, 288, 288, 288, 48, 
    288, 1, 1, 48, 288, 1, 1, 288, 96, 1, 1, 288, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 96, 96, 96, 1, 288, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 96, 232, 1, 1, 1, 1, 96, 288, 1, 1, 45, 1, 1, 96, 96, 1, 1, 1, 1, 96, 
    1, 24, 96, 96, 1, 1, 24, 1, 96, 1, 1, 24, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 
    96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 890, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1440, 1, 1, 96, 
    24, 96, 1, 1, 1, 1, 96, 96, 1, 78, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 
    1, 1, 24, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 96, 96, 96, 96, 96, 96, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 80, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 144, 144, 144, 144, 96, 144, 
    144, 144, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 10, 11, 1, 23, 1, 4, 
    1, 1, 18, 1, 18, 144, 144, 96, 1, 96, 144, 1, 1, 96 ;

 v00062_value =
  1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 91, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 20, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 48, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 86, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 48, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 23, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 56, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    92, 1, 1, 1, 1, 24, 1, 96, 96, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 
    96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1378, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 71, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 112, 1, 1, 1, 1, 1, 1, 1, 1, 1, 108, 1, 104, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 131, 1, 1, 1, 127, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 91, 
    1, 1, 1, 1, 1, 1, 1, 1, 76, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 v00054_value =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 23, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 56, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 71, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 46, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 v00060_validated =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 288, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 288, 1, 96, 1, 
    1, 288, 1, 85, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 288, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 288, 96, 1, 96, 1, 96, 1, 96, 1, 1, 86, 1, 92, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 95, 1, 1, 1, 96, 96, 1, 1, 96, 96, 
    1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 132, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 93, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 89, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 
    1, 144, 1, 1, 1, 151, 1, 1, 1, 87, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 144, 
    1, 1, 1, 111, 1, 1, 1, 144, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 73, 1, 96, 1, 1, 96, 96, 1, 95, 
    1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 144, 1, 144, 1, 1, 1, 1, 1, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 144, 1, 144, 1, 1, 1, 1, 1, 144, 1, 144, 1, 1, 1, 
    1, 1, 144, 1, 1, 1, 144, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    144, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 95, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 288, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 95, 1, 1, 96, 84, 1, 96, 1, 96, 1, 1, 96, 1, 95, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 95, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 91, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 1, 288, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 94, 1, 1, 1, 
    1, 96, 1, 1, 96, 96, 1, 288, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    288, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 288, 1, 96, 1, 96, 96, 1, 1, 1, 288, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 95, 96, 1, 96, 1, 1, 1, 96, 1, 288, 1, 96, 1, 96, 96, 1, 1, 1, 96, 
    1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 240, 1, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 288, 96, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 288, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 52, 1, 
    1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 288, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 95, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 288, 1, 1, 1, 1, 1, 40, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 288, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 288, 1, 96, 1, 288, 1, 288, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 288, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 240, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 240, 1, 96, 1, 1, 240, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 
    288, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 95, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 96, 1, 
    1, 48, 1, 1, 1, 96, 96, 1, 1, 1, 1, 48, 1, 1, 96, 1, 48, 1, 1, 1, 96, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 288, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 96, 1, 1, 96, 96, 1, 1, 92, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 53, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 240, 1, 1, 240, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 95, 1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 
    92, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 48, 1, 96, 96, 1, 1, 1, 1, 48, 1, 96, 1, 96, 1, 1, 48, 1, 1, 
    96, 48, 1, 1, 1, 1, 96, 1, 94, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 95, 95, 1, 
    1, 1, 96, 1, 96, 1, 1, 48, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 
    96, 96, 1, 1, 288, 1, 1, 1, 1, 1, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 288, 1, 1, 288, 1, 
    243, 96, 1, 96, 1, 1, 288, 96, 1, 1, 96, 288, 1, 1, 288, 1, 1439, 1, 
    1440, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 288, 1, 1, 96, 1, 
    96, 1, 96, 1, 288, 96, 1, 1, 288, 1, 166, 1, 1, 288, 1, 288, 1, 288, 288, 
    1, 1, 288, 96, 1, 1, 720, 96, 1, 1, 288, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 288, 1, 288, 96, 1, 96, 1, 95, 1, 96, 1, 1, 96, 1, 96, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 92, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 94, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 
    288, 96, 1, 96, 1, 95, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 288, 1, 288, 
    1, 288, 1, 288, 1, 288, 1, 96, 96, 1, 1, 288, 1, 1, 1, 288, 1, 1, 96, 1, 
    1, 1, 1, 288, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 288, 1, 288, 1, 
    1, 288, 1, 1, 1, 96, 1, 1, 288, 1, 1, 96, 1, 1, 288, 1, 288, 1, 96, 1, 1, 
    288, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 288, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 288, 1, 1, 96, 1, 1, 
    288, 1, 1, 95, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 288, 1, 1, 96, 288, 1, 1, 
    1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 95, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 66, 1, 1, 1, 1, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 288, 1, 288, 1, 288, 1, 96, 1, 288, 1, 1, 288, 1, 288, 1, 96, 1, 
    288, 1, 288, 1, 288, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 48, 1, 1, 48, 1, 1, 96, 24, 1, 1, 1, 96, 96, 1, 
    1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 288, 1, 288, 1, 288, 1, 288, 1, 
    96, 288, 1, 1, 288, 1, 288, 1, 288, 1, 288, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 288, 1, 1, 288, 1, 288, 288, 1, 1, 
    288, 1, 1, 288, 1, 288, 1, 1, 288, 1, 1, 288, 1, 1, 288, 1, 1, 1, 288, 1, 
    288, 1, 288, 288, 1, 288, 1, 1, 288, 1, 288, 1, 288, 1, 288, 288, 1, 1, 
    1, 1, 288, 1, 288, 1, 1, 288, 1, 288, 1, 96, 1, 288, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 24, 1, 1, 96, 1, 96, 1, 96, 1, 1, 24, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 96, 1, 96, 1, 96, 24, 
    1, 1, 1, 24, 96, 1, 1, 24, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 91, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 24, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 72, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 95, 1, 1, 95, 1, 96, 1, 1, 95, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 94, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 94, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 24, 
    96, 1, 96, 1, 1, 48, 24, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 1, 1, 1, 95, 94, 1, 1, 96, 96, 1, 96, 1, 1, 83, 1, 1, 96, 1, 
    48, 1, 48, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 48, 1, 24, 1, 24, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 24, 1, 1, 1, 1, 48, 96, 1, 1, 1, 24, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    24, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    24, 1, 48, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 288, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 48, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 24, 1, 1, 48, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 221, 1, 1, 96, 1, 89, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 264, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 
    1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 95, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 84, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 96, 24, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 96, 1, 1, 1, 1, 1, 87, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 203, 1, 1, 1, 1, 1, 1, 1, 24, 1, 24, 1, 24, 1, 92, 1, 24, 
    1, 24, 1, 1, 95, 96, 1, 1, 96, 96, 1, 96, 1, 1, 24, 48, 1, 48, 1, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 24, 1, 24, 1, 1, 24, 1, 
    96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 
    92, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 24, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 24, 1, 1, 24, 24, 1, 1, 1, 1, 24, 1, 96, 1, 24, 1, 96, 1, 1, 
    96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 24, 1, 1, 24, 1, 23, 1, 24, 1, 
    1, 24, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 24, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 24, 1, 1, 24, 1, 24, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 91, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 95, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 92, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 93, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 24, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 94, 1, 1, 92, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 48, 24, 
    1, 1, 96, 1, 1, 48, 48, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 48, 1, 24, 1, 1, 
    96, 1, 1, 1, 24, 1, 1, 48, 24, 1, 1, 48, 48, 1, 96, 1, 1, 96, 1, 96, 48, 
    1, 48, 1, 96, 1, 48, 1, 96, 1, 1, 96, 1, 48, 1, 48, 1, 96, 1, 24, 1, 48, 
    1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 48, 1, 1, 48, 1, 48, 96, 1, 96, 
    1, 1, 1, 48, 1, 48, 1, 96, 1, 24, 1, 1, 48, 1, 1, 96, 1, 48, 48, 1, 1, 
    96, 1, 1, 56, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 95, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 95, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 48, 1, 48, 1, 1, 48, 
    1, 1, 1, 1, 96, 48, 1, 48, 1, 1, 48, 1, 48, 1, 48, 1, 1, 48, 1, 1, 96, 
    96, 1, 1, 96, 1, 1, 1, 48, 1, 1, 1, 48, 48, 1, 95, 1, 1, 1, 96, 1, 48, 1, 
    48, 1, 48, 1, 47, 1, 1, 96, 1, 96, 24, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 
    48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 44, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 24, 1, 1, 48, 
    1, 1, 24, 1, 1, 1, 1, 96, 24, 1, 1, 1, 96, 1, 96, 1, 96, 1, 24, 1, 1, 96, 
    96, 1, 1, 1, 96, 1, 80, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 24, 1, 1, 24, 
    1, 96, 1, 1, 1, 96, 24, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 48, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 288, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 96, 1, 96, 1, 1, 90, 1, 1, 48, 1, 1, 24, 1, 1, 48, 1, 1, 1, 48, 1, 
    96, 1, 48, 1, 96, 1, 48, 1, 93, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 25, 1, 96, 1, 93, 1, 1, 1, 95, 1, 96, 1, 82, 1, 96, 1, 1, 81, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 24, 1, 1, 48, 1, 48, 1, 48, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 91, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 95, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 89, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    24, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 48, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 48, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 93, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 48, 1, 1, 95, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 95, 1, 1, 96, 1, 95, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 84, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 288, 1, 96, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 48, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 24, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 
    1, 1, 95, 1, 1, 1, 1, 96, 96, 1, 1, 48, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 1, 1, 48, 1, 48, 1, 96, 1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 96, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 96, 
    1, 1, 48, 1, 1, 1, 96, 1, 48, 1, 1, 24, 48, 1, 1, 96, 1, 1, 1, 48, 1, 96, 
    1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 96, 1, 1, 48, 1, 63, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 96, 1, 1, 96, 1, 1, 1, 48, 1, 
    96, 1, 1, 1, 96, 1, 48, 1, 48, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 48, 
    1, 1, 48, 1, 1, 96, 1, 1, 96, 1, 1, 1, 48, 1, 1, 96, 1, 48, 1, 1, 96, 1, 
    1, 95, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 48, 48, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 48, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 48, 1, 1, 1, 1, 46, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 1, 42, 1, 1, 
    1, 48, 1, 1, 47, 1, 1, 1, 47, 1, 1, 1, 96, 1, 48, 1, 48, 48, 1, 1, 1, 1, 
    96, 1, 1, 1, 48, 1, 48, 1, 48, 1, 1, 1, 48, 1, 48, 1, 96, 1, 48, 1, 1, 
    96, 1, 48, 48, 1, 1, 48, 1, 1, 1, 48, 1, 47, 1, 1, 1, 1, 48, 46, 1, 1, 
    96, 1, 48, 24, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 48, 1, 1, 1, 96, 96, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 
    1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 288, 1, 1, 288, 1, 1, 264, 1, 1, 96, 1, 
    1, 95, 1, 1, 92, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 288, 1, 1, 
    288, 1, 1, 96, 1, 96, 1, 288, 1, 1, 288, 288, 1, 1, 1, 288, 1, 1, 1, 288, 
    1, 288, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 144, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 93, 1, 1, 1, 96, 1, 1, 92, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    95, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 92, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 1, 90, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 95, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 95, 96, 1, 1, 1, 1, 1, 1, 1, 48, 1, 
    48, 1, 1, 1, 48, 96, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 48, 1, 1, 
    1, 48, 1, 1, 48, 92, 1, 96, 1, 1, 1, 48, 1, 1, 1, 96, 1, 1, 1, 96, 48, 1, 
    1, 1, 1, 1, 48, 1, 1, 91, 1, 48, 1, 1, 1, 1, 1, 48, 1, 48, 1, 1, 1, 48, 
    48, 1, 1, 1, 1, 1, 97, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 97, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 94, 1, 1, 1, 1, 
    1, 1, 97, 1, 1, 97, 1, 1, 96, 1, 48, 1, 96, 1, 1, 96, 96, 1, 1, 48, 1, 1, 
    43, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 48, 1, 1, 1, 1, 48, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 48, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 48, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 48, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 48, 1, 95, 1, 1, 96, 1, 96, 
    96, 1, 48, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 
    1, 1, 48, 1, 96, 1, 1, 96, 1, 48, 1, 1, 1, 96, 96, 1, 1, 95, 1, 1, 288, 
    1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 93, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 24, 1, 1, 96, 96, 1, 1, 22, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 24, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 
    96, 1, 1, 94, 1, 96, 1, 96, 1, 1, 96, 1, 1, 24, 1, 96, 24, 1, 1, 96, 1, 
    96, 96, 1, 1, 1, 96, 1, 24, 49, 1, 1, 96, 1, 96, 1, 1, 1, 1, 48, 1, 1, 
    288, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 9, 1, 1, 1, 96, 1, 288, 
    1, 288, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 24, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 288, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 288, 1, 1, 96, 1, 1, 288, 1, 1, 1, 96, 1, 135, 1, 96, 
    1, 1, 1, 288, 1, 1, 96, 1, 1, 34, 1, 1, 95, 1, 1, 96, 1, 1, 288, 96, 1, 
    96, 1, 1, 1, 93, 1, 1, 1, 96, 1, 1, 288, 1, 1, 1, 288, 1, 1, 96, 1, 1, 1, 
    1, 288, 1, 1, 288, 1, 1, 288, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 264, 287, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 288, 1, 1, 96, 1, 1, 273, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 48, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 120, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 92, 1, 96, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 120, 
    1, 1, 1, 120, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 45, 1, 1, 240, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 288, 96, 1, 1, 96, 96, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 48, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 
    96, 1, 1, 48, 1, 1, 48, 1, 97, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 48, 96, 1, 1, 96, 1, 
    93, 1, 1, 48, 1, 48, 1, 1, 48, 1, 48, 48, 1, 96, 1, 1, 48, 1, 96, 96, 1, 
    1, 1, 48, 1, 96, 1, 96, 1, 48, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 288, 1, 
    1, 96, 1, 48, 1, 96, 1, 96, 1, 96, 1, 288, 1, 96, 1, 96, 1, 288, 96, 1, 
    1, 1, 1, 48, 1, 1, 96, 1, 1, 144, 1, 96, 1, 1, 1, 48, 1, 48, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 99, 1, 99, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 97, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 98, 1, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 1, 288, 1, 288, 96, 1, 94, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 81, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 26, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 10, 1, 
    96, 1, 95, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 89, 1, 1, 96, 
    1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 48, 1, 48, 1, 96, 1, 96, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 74, 1, 96, 1, 96, 1, 48, 96, 
    1, 48, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 25, 1, 1, 1, 96, 1, 88, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 47, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 82, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 14, 1, 1, 96, 1, 
    24, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 95, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    288, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 88, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 87, 57, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 144, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    288, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 288, 1, 96, 96, 1, 96, 1, 96, 1, 
    288, 1, 1, 1, 288, 96, 1, 1, 1, 1, 1, 288, 1, 96, 1, 1, 1, 288, 1, 1, 96, 
    1, 1, 1, 1, 189, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 144, 
    1, 1, 1, 96, 1, 1, 1, 288, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 90, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 81, 1, 96, 1, 96, 1, 96, 1, 1, 82, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 86, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 13, 90, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 92, 1, 96, 1, 1, 1, 96, 96, 1, 1, 8, 96, 1, 
    96, 1, 96, 1, 144, 1, 96, 1, 58, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 48, 48, 1, 1, 96, 1, 1, 47, 
    46, 1, 1, 1, 48, 1, 48, 1, 48, 1, 48, 1, 48, 1, 1, 1, 1, 48, 1, 1, 48, 
    96, 1, 48, 1, 1, 1, 288, 1, 1, 288, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 95, 1, 95, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 1, 96, 96, 1, 95, 1, 1, 1, 288, 1, 1, 1, 96, 1, 1, 288, 1, 1, 1, 
    1, 288, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 95, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 144, 1, 144, 1, 1, 1, 96, 1, 48, 1, 1, 96, 1, 1, 288, 1, 
    278, 1, 1, 96, 1, 96, 1, 1, 288, 1, 288, 1, 288, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 288, 1, 96, 
    1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 288, 1, 288, 1, 1, 
    1, 75, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 24, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 286, 1, 1, 96, 1, 1, 96, 96, 1, 1, 93, 1, 
    96, 1, 96, 1, 94, 48, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 95, 1, 96, 1, 96, 95, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 94, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 
    1, 1, 69, 1, 49, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 58, 
    96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 95, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 61, 1, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 34, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 35, 1, 1, 86, 1, 96, 
    1, 1, 96, 96, 1, 96, 1, 95, 1, 96, 1, 1, 88, 1, 96, 96, 1, 1, 96, 1, 96, 
    94, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 50, 1, 1, 96, 96, 1, 
    96, 1, 73, 1, 1, 96, 57, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 95, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 37, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 95, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 92, 1, 84, 1, 32, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 288, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 288, 1, 1, 288, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 88, 1, 96, 1, 96, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 288, 1, 288, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 95, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 62, 
    1, 96, 89, 1, 96, 1, 1, 96, 1, 1, 1, 1, 92, 1, 96, 1, 1, 1, 1, 96, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 87, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 95, 1, 1, 1, 
    1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 70, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 14, 1, 1, 1, 96, 1, 96, 1, 1, 49, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 25, 1, 1, 96, 
    1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 33, 1, 1, 97, 1, 
    1, 1, 1, 1, 1, 93, 1, 1, 1, 1, 89, 1, 1, 88, 1, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 88, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 
    1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 96, 1, 288, 1, 1, 288, 1, 288, 96, 
    1, 1, 1, 288, 1, 288, 1, 1, 288, 1, 288, 1, 288, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 288, 1, 42, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 288, 
    1, 288, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 288, 1, 1, 172, 1, 96, 96, 1, 
    1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    29, 1, 1, 94, 96, 1, 1, 89, 96, 1, 1, 96, 95, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 95, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 90, 1, 96, 1, 1, 71, 1, 
    95, 96, 1, 1, 1, 96, 1, 96, 1, 52, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 
    1, 49, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 288, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 
    1, 96, 1, 94, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 95, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 81, 1, 96, 96, 1, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 88, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 90, 1, 1, 
    288, 1, 1, 4, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 94, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 89, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 92, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 69, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 54, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 36, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 94, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 97, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 94, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 288, 1, 288, 1, 1, 288, 
    1, 264, 92, 1, 1, 1, 288, 96, 1, 1, 1, 288, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 288, 1, 1, 288, 1, 288, 288, 1, 1, 1, 288, 1, 
    288, 1, 24, 1, 1, 1, 1, 1, 281, 1, 288, 288, 1, 1, 1, 287, 1, 288, 1, 
    288, 1, 288, 1, 1, 24, 288, 1, 1, 285, 1, 288, 1, 1, 264, 1, 288, 1, 288, 
    1, 288, 288, 1, 1, 288, 1, 1, 264, 1, 290, 288, 1, 1, 288, 288, 1, 1, 96, 
    1, 1, 1, 48, 1, 96, 1, 1, 1, 48, 96, 1, 1, 1, 47, 1, 96, 1, 1, 1, 48, 94, 
    1, 1, 1, 48, 264, 1, 1, 288, 1, 1, 1, 288, 1, 288, 288, 1, 1, 1, 288, 
    255, 1, 1, 287, 1, 48, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 46, 1, 96, 1, 1, 
    94, 96, 1, 24, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 48, 
    1, 1, 24, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 1, 48, 1, 24, 1, 48, 1, 1, 1, 24, 
    96, 1, 1, 1, 1, 277, 89, 1, 24, 1, 1, 1, 288, 1, 1, 288, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 288, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    22, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 95, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 98, 1, 1, 96, 
    47, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 92, 1, 1, 55, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 
    1, 1, 1, 96, 24, 1, 1, 96, 1, 1, 1, 24, 1, 1, 286, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 156, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 85, 1, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 86, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 
    1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 48, 1, 1, 96, 1, 48, 1, 1, 24, 48, 1, 1, 1, 96, 1, 
    1, 1, 48, 1, 96, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 96, 48, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 24, 1, 1, 48, 1, 1, 96, 1, 92, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 24, 1, 1, 1, 96, 1, 96, 96, 
    1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 48, 1, 96, 1, 1, 48, 1, 1, 96, 1, 1, 26, 
    1, 1, 1, 1, 96, 1, 96, 1, 48, 1, 48, 1, 1, 1, 1, 1, 48, 24, 1, 1, 95, 1, 
    96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 70, 1, 48, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 48, 1, 1, 24, 1, 1, 1, 
    96, 92, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 94, 1, 96, 1, 1, 
    24, 96, 1, 48, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 48, 1, 1, 96, 1, 1, 94, 1, 1, 48, 1, 1, 96, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 96, 
    1, 1, 1, 288, 1, 96, 1, 1, 1, 1, 290, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 24, 1, 96, 1, 1, 96, 1, 1, 96, 1, 48, 1, 1, 96, 1, 1, 24, 1, 1, 
    96, 1, 48, 1, 1, 96, 1, 1, 1, 1, 1, 48, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 92, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 48, 1, 1, 48, 48, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 1, 96, 48, 1, 1, 1, 1, 48, 96, 1, 
    1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 24, 
    1, 48, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 
    48, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 48, 1, 1, 1, 
    48, 1, 96, 1, 1, 48, 1, 1, 1, 96, 1, 48, 1, 48, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 93, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 70, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 1, 1, 
    30, 1, 24, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    15, 1, 1, 96, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 86, 1, 1, 60, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 
    1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    96, 1, 48, 1, 1, 48, 1, 1, 1, 48, 1, 48, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    62, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 93, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 48, 1, 37, 1, 1, 1, 48, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 48, 1, 48, 1, 1, 96, 1, 1, 95, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 48, 1, 1, 96, 1, 96, 1, 96, 48, 1, 1, 1, 96, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 144, 1, 24, 1, 1, 1, 1, 96, 24, 1, 1, 1, 
    48, 1, 1, 1, 96, 1, 1, 48, 1, 24, 1, 96, 1, 1, 46, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 24, 96, 96, 1, 1, 1, 1, 24, 1, 
    1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 24, 1, 1, 48, 1, 24, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 90, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 48, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 285, 1, 1, 1, 288, 1, 288, 1, 1, 96, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 24, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 95, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 96, 48, 1, 1, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 48, 1, 1, 48, 1, 1, 48, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 48, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 56, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 48, 1, 1, 48, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 
    1, 1, 1, 1, 1, 40, 48, 1, 1, 48, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 48, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 96, 1, 1, 95, 96, 1, 1, 96, 1, 85, 1, 1, 1, 48, 1, 96, 
    1, 1, 1, 1, 92, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 88, 96, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 95, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 73, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    94, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 94, 96, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 95, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 95, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 87, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 6, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 26, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 60, 1, 1, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 90, 1, 1, 96, 1, 96, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 95, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 95, 1, 1, 288, 1, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 288, 1, 1, 95, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    288, 1, 96, 1, 1, 1, 96, 1, 288, 1, 1, 1, 288, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 288, 1, 1, 288, 95, 
    1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 95, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 288, 
    1, 288, 1, 1, 1, 96, 1, 1, 288, 1, 1, 288, 1, 1, 96, 1, 1, 1, 288, 1, 1, 
    288, 1, 1, 96, 1, 288, 1, 288, 1, 288, 1, 288, 1, 288, 1, 288, 1, 288, 1, 
    288, 1, 1, 288, 96, 1, 1, 1, 1, 288, 1, 288, 288, 1, 1, 288, 1, 288, 288, 
    1, 1, 288, 1, 288, 1, 1, 1, 1, 1, 288, 1, 288, 1, 288, 1, 1, 1, 288, 196, 
    1, 1, 288, 288, 1, 1, 288, 288, 1, 1, 288, 288, 1, 288, 1, 288, 1, 288, 
    1, 288, 1, 1, 288, 1, 1, 96, 288, 1, 1, 1, 288, 1, 1, 1, 1, 96, 1, 1, 96, 
    96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 93, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 95, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 68, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 92, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 95, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 11, 
    1, 1, 96, 288, 1, 1, 1, 96, 1, 1, 96, 96, 1, 288, 1, 288, 1, 1, 1, 96, 1, 
    96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 93, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 
    16, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 144, 1, 
    1, 1, 288, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 95, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 96, 64, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 80, 
    96, 1, 1, 4, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 1, 93, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 93, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 288, 1, 1, 96, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 
    96, 1, 1, 96, 94, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 92, 1, 1, 94, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 90, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 91, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 94, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 101, 1, 1, 1, 
    93, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 94, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 96, 1, 1, 94, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 
    1, 1, 1, 96, 96, 1, 96, 1, 95, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 95, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 192, 
    1, 1, 96, 1, 192, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 81, 1, 96, 1, 
    44, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 65, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 53, 1, 1, 1, 1, 96, 1, 95, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 98, 1, 96, 1, 1, 96, 1, 1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 95, 1, 1, 1, 1, 164, 1, 96, 1, 96, 1, 96, 97, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 100, 1, 96, 96, 1, 99, 1, 96, 1, 1, 96, 96, 1, 1, 97, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 97, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    94, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 62, 96, 1, 1, 96, 96, 96, 96, 96, 96, 
    96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 94, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 92, 1, 90, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 92, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 35, 1, 1, 1, 1, 
    43, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 76, 1, 1, 1, 1, 1, 96, 96, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 80, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 15, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 95, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 89, 1, 96, 1, 76, 1, 96, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 85, 1, 96, 1, 96, 1, 96, 1, 62, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 90, 1, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 95, 1, 96, 1, 1, 95, 1, 1, 1, 98, 1, 96, 
    1, 100, 1, 96, 1, 96, 1, 96, 1, 1, 96, 98, 1, 1, 96, 1, 96, 96, 1, 96, 1, 
    96, 1, 94, 1, 32, 1, 288, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 
    1, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 93, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 49, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 96, 1, 96, 1, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    94, 1, 1, 95, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 85, 1, 85, 1, 85, 1, 85, 1, 1, 85, 86, 1, 
    82, 82, 1, 82, 1, 1, 82, 82, 1, 1, 1, 82, 1, 82, 1, 82, 1, 86, 1, 96, 1, 
    96, 1, 1, 96, 86, 1, 86, 1, 86, 1, 86, 87, 1, 59, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 93, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 84, 1, 1, 1, 84, 1, 84, 1, 78, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 96, 96, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 35, 
    1, 1, 96, 1, 96, 1, 1, 1, 84, 1, 84, 1, 1, 1, 1, 84, 84, 1, 1, 1, 84, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 84, 1, 1, 89, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 54, 1, 1, 96, 1, 96, 1, 83, 1, 1, 
    1, 75, 1, 1, 1, 1, 96, 1, 96, 1, 1, 72, 96, 1, 1, 1, 96, 96, 1, 1, 20, 
    96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    60, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 144, 1, 48, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 227, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 144, 1, 144, 1, 144, 1, 144, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 91, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 53, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 32, 1, 86, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 24, 1, 96, 1, 24, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 48, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 95, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 94, 1, 96, 1, 
    66, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 93, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 56, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 288, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 97, 
    1, 96, 95, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 19, 1, 1, 
    96, 1, 96, 1, 96, 1, 43, 1, 11, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 83, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 89, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 97, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 56, 1, 1, 84, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 99, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 41, 1, 96, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 52, 1, 96, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 28, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 44, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 86, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 48, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 89, 1, 
    1, 1, 48, 1, 1, 48, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 98, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 97, 1, 1, 96, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 114, 1, 1, 108, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    106, 1, 96, 1, 1, 1, 96, 1, 1, 112, 1, 1, 1, 1, 107, 1, 1, 1, 1, 1, 1, 1, 
    137, 1, 1, 126, 1, 128, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 94, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 288, 1, 1, 97, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 95, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 1, 48, 1, 96, 1, 1, 42, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 87, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 88, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 15, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 64, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 94, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 225, 96, 1, 96, 1, 96, 1, 96, 1, 
    112, 1, 96, 1, 102, 1, 100, 1, 96, 1, 96, 1, 288, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 52, 96, 1, 1, 1, 1, 14, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 84, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 58, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 137, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 88, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 288, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 890, 1, 1, 96, 1, 1, 96, 1, 89, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 288, 1, 1193, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 88, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1 ;

 v00065_validated =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 96, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 288, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 288, 1, 1, 1, 96, 
    288, 1, 85, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 96, 1, 
    96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 288, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 288, 1, 1, 96, 1, 96, 1, 96, 1, 96, 86, 1, 92, 
    1, 1, 96, 1, 96, 96, 1, 92, 96, 1, 96, 1, 1, 95, 96, 96, 1, 1, 96, 96, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 144, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 93, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 89, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 96, 1, 1, 96, 
    1, 96, 144, 1, 1, 1, 151, 1, 1, 1, 87, 1, 1, 1, 97, 1, 1, 1, 1, 1, 1, 1, 
    144, 1, 1, 1, 111, 1, 1, 1, 144, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 73, 1, 96, 96, 1, 
    1, 96, 1, 95, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 
    144, 1, 1, 96, 1, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 144, 
    1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 144, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 95, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 95, 96, 1, 1, 84, 1, 96, 1, 96, 96, 1, 95, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 91, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 288, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 288, 1, 1, 
    1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 94, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 288, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 288, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 96, 1, 96, 1, 96, 96, 1, 48, 45, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 96, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    72, 1, 96, 96, 1, 1, 96, 96, 1, 96, 96, 96, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 96, 1, 288, 1, 96, 1, 96, 1, 1, 96, 
    96, 288, 1, 12, 1, 96, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 
    288, 288, 1, 288, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 95, 1, 1, 96, 1, 
    96, 1, 96, 1, 288, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 96, 1, 1, 96, 240, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 288, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 288, 96, 1, 96, 1, 1, 96, 1, 96, 96, 52, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 288, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 95, 1, 96, 1, 96, 1, 96, 96, 
    96, 1, 96, 1, 1, 288, 1, 1, 288, 1, 1, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 96, 288, 1, 288, 288, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 288, 1, 288, 240, 1, 1, 288, 288, 1, 96, 1, 96, 1, 96, 96, 1, 
    1, 96, 96, 96, 1, 1, 288, 1, 96, 1, 288, 1, 288, 1, 1, 96, 1, 96, 96, 1, 
    96, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 96, 96, 1, 96, 96, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 288, 
    96, 1, 96, 1, 96, 96, 96, 96, 1, 96, 1, 1, 96, 96, 1, 119, 1, 240, 1, 1, 
    96, 1, 96, 185, 1, 1, 96, 1, 96, 240, 1, 1, 96, 96, 1, 1, 1, 240, 1, 1, 
    96, 240, 1, 240, 1, 1, 1, 96, 96, 1, 240, 1, 1, 240, 1, 1, 1, 96, 240, 1, 
    1, 240, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 240, 1, 240, 1, 230, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 96, 240, 1, 240, 1, 237, 1, 240, 1, 240, 1, 
    240, 1, 240, 1, 96, 1, 1, 96, 240, 1, 96, 206, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 
    1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 288, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 
    96, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 96, 96, 1, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 95, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 1, 
    96, 1, 1, 48, 1, 96, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 96, 1, 48, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 288, 1, 96, 96, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 92, 1, 240, 1, 1, 239, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 53, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 240, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 96, 240, 1, 1, 1, 1, 1, 1, 240, 1, 96, 1, 96, 1, 1, 240, 240, 1, 
    1, 240, 96, 1, 240, 240, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 
    240, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 
    1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 95, 
    1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 
    1, 96, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 96, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 92, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 48, 1, 96, 1, 1, 96, 1, 1, 
    48, 1, 96, 1, 96, 1, 1, 48, 1, 1, 96, 1, 1, 48, 1, 1, 96, 1, 94, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 95, 1, 1, 95, 1, 1, 1, 96, 1, 96, 48, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    1, 1, 96, 96, 1, 240, 240, 96, 1, 1, 96, 96, 1, 1, 96, 288, 1, 1, 1, 1, 
    1, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 288, 288, 1, 243, 1, 1, 96, 1, 96, 288, 1, 1, 
    96, 96, 1, 1, 288, 288, 1, 1439, 1, 1440, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 96, 1, 1, 288, 96, 1, 96, 1, 96, 1, 288, 1, 1, 96, 288, 1, 
    166, 1, 288, 288, 1, 288, 1, 288, 1, 1, 288, 288, 1, 1, 96, 720, 1, 1, 
    96, 288, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 288, 1, 288, 1, 1, 96, 
    1, 96, 1, 95, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 288, 1, 96, 96, 1, 96, 96, 1, 
    1, 96, 1, 96, 1, 96, 96, 1, 92, 1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 94, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 288, 1, 1, 96, 1, 96, 1, 
    95, 96, 1, 1, 96, 1, 96, 96, 1, 96, 288, 1, 288, 1, 288, 1, 288, 1, 288, 
    1, 96, 1, 1, 96, 288, 1, 1, 1, 288, 1, 1, 1, 1, 96, 1, 1, 288, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 288, 1, 288, 1, 288, 1, 1, 1, 1, 288, 1, 1, 1, 
    96, 288, 1, 1, 1, 1, 96, 1, 1, 288, 1, 288, 1, 96, 288, 1, 1, 1, 1, 96, 
    265, 1, 1, 1, 96, 288, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 288, 1, 1, 288, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 
    96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 96, 1, 1, 
    1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 288, 1, 1, 1, 1, 
    96, 288, 1, 1, 95, 1, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 288, 1, 1, 96, 1, 1, 
    1, 288, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 96, 1, 1, 95, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 66, 
    1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 96, 288, 1, 288, 1, 288, 1, 96, 1, 288, 1, 288, 
    288, 1, 288, 1, 96, 1, 288, 1, 288, 1, 288, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 48, 48, 1, 96, 1, 
    1, 1, 24, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 288, 1, 
    288, 1, 288, 1, 288, 1, 96, 1, 1, 288, 288, 1, 288, 1, 288, 1, 288, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 288, 
    288, 1, 288, 1, 1, 288, 288, 1, 288, 288, 1, 288, 1, 288, 288, 1, 288, 
    288, 1, 288, 288, 1, 288, 288, 288, 1, 288, 1, 288, 1, 1, 288, 1, 288, 
    288, 1, 288, 1, 288, 1, 288, 1, 1, 288, 288, 288, 288, 1, 288, 1, 288, 
    288, 1, 288, 1, 96, 1, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 
    1, 1, 1, 24, 96, 1, 96, 1, 96, 1, 1, 1, 1, 24, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 24, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 96, 96, 96, 96, 96, 1, 96, 96, 24, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 96, 96, 93, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 96, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    96, 96, 1, 1, 96, 96, 96, 1, 1, 96, 1, 1, 1, 96, 24, 1, 96, 1, 96, 1, 96, 
    1, 1, 24, 1, 24, 1, 1, 96, 24, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 95, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 91, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 24, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 72, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 95, 1, 1, 96, 1, 1, 95, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 94, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 94, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 73, 
    1, 1, 1, 96, 96, 1, 24, 1, 1, 96, 1, 96, 48, 1, 1, 24, 1, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 95, 1, 1, 94, 96, 1, 1, 96, 
    1, 96, 84, 1, 1, 1, 1, 96, 1, 48, 1, 48, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 48, 1, 24, 1, 24, 1, 24, 24, 1, 96, 96, 24, 24, 24, 24, 96, 96, 
    1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 24, 1, 24, 24, 48, 48, 1, 1, 96, 24, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 24, 1, 24, 96, 1, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 24, 1, 48, 96, 96, 1, 1, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 24, 24, 1, 96, 96, 1, 
    96, 1, 48, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 24, 1, 
    1, 48, 1, 1, 24, 24, 1, 24, 48, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 221, 92, 1, 96, 1, 89, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 24, 24, 96, 96, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    264, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 95, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 95, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 96, 
    1, 95, 94, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 96, 96, 96, 1, 
    96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 203, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 24, 1, 24, 1, 24, 1, 92, 1, 24, 1, 24, 95, 1, 1, 96, 96, 1, 1, 96, 1, 
    96, 24, 1, 1, 48, 1, 48, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 96, 1, 96, 96, 96, 1, 96, 96, 1, 96, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 1, 24, 1, 24, 24, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 24, 96, 1, 1, 96, 1, 92, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 24, 96, 1, 96, 1, 1, 1, 96, 1, 1, 24, 24, 1, 1, 24, 96, 
    1, 1, 1, 24, 1, 96, 1, 24, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 96, 1, 1, 1, 1, 1, 
    1, 24, 1, 24, 24, 1, 24, 1, 23, 1, 24, 24, 1, 96, 1, 24, 96, 96, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 24, 96, 1, 1, 1, 96, 1, 1, 24, 1, 1, 96, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 24, 24, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 91, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 95, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 95, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 92, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 93, 1, 1, 96, 1, 96, 1, 1, 1, 1, 92, 1, 96, 1, 1, 
    24, 1, 96, 1, 96, 1, 24, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 94, 1, 1, 92, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 48, 1, 1, 24, 1, 1, 
    96, 48, 1, 1, 48, 1, 24, 1, 1, 1, 96, 1, 1, 23, 1, 48, 1, 24, 24, 1, 96, 
    1, 1, 1, 24, 48, 1, 1, 24, 48, 1, 1, 48, 1, 96, 96, 1, 96, 1, 1, 48, 1, 
    48, 1, 96, 1, 48, 1, 96, 96, 1, 1, 1, 48, 1, 48, 1, 96, 1, 24, 1, 48, 96, 
    1, 96, 1, 1, 96, 96, 1, 1, 96, 48, 1, 1, 48, 1, 48, 1, 1, 96, 1, 96, 1, 
    48, 1, 48, 1, 96, 1, 24, 1, 96, 48, 1, 48, 96, 1, 48, 1, 1, 48, 1, 1, 96, 
    1, 1, 56, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 
    95, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 95, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 48, 1, 48, 48, 1, 
    48, 48, 48, 96, 1, 1, 48, 1, 48, 48, 1, 48, 1, 48, 1, 48, 1, 1, 48, 96, 
    1, 1, 96, 96, 1, 1, 48, 48, 1, 48, 48, 48, 1, 1, 48, 1, 95, 1, 96, 1, 1, 
    1, 48, 1, 48, 1, 48, 1, 47, 96, 1, 96, 1, 1, 24, 48, 48, 1, 1, 1, 24, 1, 
    48, 96, 1, 48, 24, 1, 24, 1, 48, 24, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 
    1, 24, 24, 1, 48, 24, 1, 24, 1, 24, 96, 1, 1, 24, 24, 96, 1, 96, 1, 96, 
    1, 24, 1, 1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 24, 24, 1, 96, 96, 1, 96, 
    24, 24, 96, 1, 1, 24, 24, 1, 24, 1, 96, 96, 96, 1, 1, 24, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 1, 48, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 288, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 96, 
    1, 1, 96, 96, 1, 24, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 96, 1, 90, 94, 1, 
    48, 96, 1, 23, 24, 1, 48, 24, 48, 1, 96, 1, 24, 1, 48, 1, 48, 1, 93, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 25, 1, 96, 1, 93, 1, 1, 1, 
    95, 1, 96, 1, 82, 1, 96, 1, 96, 81, 1, 96, 96, 1, 96, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 24, 48, 1, 48, 1, 48, 1, 96, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 91, 1, 1, 96, 96, 96, 96, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 95, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 96, 96, 96, 96, 1, 1, 96, 2, 96, 1, 1, 96, 96, 96, 1, 96, 1, 1, 96, 
    1, 96, 89, 1, 1, 1, 48, 1, 1, 1, 96, 96, 1, 96, 96, 1, 1, 48, 1, 1, 48, 
    1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 76, 36, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 24, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 48, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 96, 96, 1, 96, 1, 1, 1, 48, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 93, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 
    96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 95, 96, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 94, 95, 92, 96, 96, 1, 96, 96, 96, 1, 1, 96, 48, 48, 48, 96, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 48, 1, 1, 
    95, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 96, 48, 48, 1, 1, 96, 96, 96, 1, 
    95, 1, 1, 96, 1, 1, 1, 95, 48, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 48, 1, 84, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 96, 1, 1, 1, 96, 96, 
    96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 288, 1, 96, 1, 1, 96, 1, 
    1, 96, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 288, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 96, 94, 1, 96, 
    96, 96, 1, 1, 85, 88, 1, 96, 1, 96, 48, 1, 48, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 48, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 48, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 94, 
    1, 24, 96, 1, 42, 43, 1, 1, 96, 288, 1, 96, 1, 44, 40, 1, 96, 1, 1, 288, 
    1, 1, 96, 96, 1, 1, 96, 1, 96, 95, 1, 47, 48, 1, 96, 1, 1, 96, 48, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 48, 1, 48, 1, 96, 1, 48, 1, 48, 1, 
    48, 96, 1, 1, 48, 48, 1, 48, 48, 1, 95, 48, 89, 48, 48, 48, 48, 1, 96, 1, 
    48, 48, 48, 48, 48, 1, 48, 48, 1, 48, 1, 96, 48, 1, 48, 48, 96, 1, 48, 1, 
    48, 24, 1, 1, 48, 96, 1, 1, 96, 48, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 48, 1, 48, 48, 1, 96, 48, 1, 63, 1, 96, 1, 48, 1, 1, 96, 1, 96, 
    48, 48, 1, 48, 1, 48, 1, 48, 1, 96, 96, 1, 96, 1, 48, 1, 96, 1, 48, 48, 
    96, 1, 48, 1, 48, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 69, 1, 48, 1, 
    1, 48, 33, 1, 96, 96, 1, 1, 1, 96, 1, 48, 96, 1, 96, 1, 48, 1, 1, 96, 96, 
    1, 95, 96, 1, 1, 1, 96, 1, 48, 1, 1, 96, 1, 1, 96, 48, 1, 1, 48, 1, 96, 
    1, 48, 1, 93, 1, 48, 1, 96, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 96, 96, 1, 96, 96, 1, 48, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 96, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 48, 1, 20, 1, 96, 1, 96, 1, 96, 
    48, 1, 48, 1, 1, 48, 48, 1, 1, 48, 1, 48, 46, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 48, 48, 1, 47, 48, 48, 1, 1, 40, 48, 1, 1, 48, 
    48, 1, 96, 48, 42, 1, 1, 1, 48, 1, 1, 47, 1, 1, 1, 47, 1, 96, 48, 96, 1, 
    48, 1, 48, 1, 1, 48, 1, 1, 96, 1, 1, 1, 48, 1, 48, 1, 48, 1, 1, 48, 48, 
    1, 48, 1, 96, 1, 48, 1, 1, 96, 1, 48, 1, 1, 48, 48, 1, 48, 48, 48, 1, 47, 
    1, 48, 48, 1, 48, 1, 1, 46, 96, 1, 48, 1, 1, 24, 96, 1, 1, 96, 1, 48, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 48, 1, 48, 24, 1, 96, 1, 96, 
    1, 1, 96, 24, 1, 96, 1, 96, 1, 288, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 97, 96, 1, 96, 1, 48, 1, 96, 
    92, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 48, 1, 96, 1, 1, 96, 95, 96, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 288, 1, 
    1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 288, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 288, 1, 1, 288, 1, 1, 264, 1, 1, 96, 1, 95, 1, 1, 1, 92, 
    1, 96, 1, 1, 96, 1, 96, 96, 96, 1, 1, 1, 96, 1, 288, 1, 1, 288, 1, 1, 96, 
    1, 96, 1, 288, 1, 1, 288, 1, 1, 288, 1, 288, 1, 1, 1, 288, 1, 1, 1, 288, 
    1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    96, 144, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 288, 1, 1, 93, 1, 96, 1, 1, 1, 1, 92, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 96, 1, 1, 
    96, 96, 1, 1, 96, 288, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 288, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 96, 288, 1, 1, 96, 1, 96, 96, 96, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 95, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 96, 96, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 
    96, 24, 24, 24, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 92, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 
    24, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 24, 24, 1, 
    90, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 
    96, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 95, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 
    96, 1, 96, 1, 96, 96, 1, 96, 95, 1, 1, 96, 96, 1, 95, 95, 48, 1, 1, 48, 
    1, 1, 48, 1, 1, 1, 96, 1, 1, 48, 1, 48, 1, 1, 48, 48, 1, 1, 48, 1, 48, 1, 
    48, 1, 48, 1, 1, 1, 92, 1, 96, 1, 1, 1, 48, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    48, 48, 1, 1, 1, 48, 1, 1, 91, 1, 48, 48, 1, 1, 48, 1, 1, 1, 48, 1, 48, 
    1, 1, 48, 1, 288, 1, 97, 1, 95, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 96, 1, 
    96, 96, 287, 1, 1, 48, 1, 96, 1, 97, 1, 1, 1, 1, 1, 96, 288, 1, 1, 288, 
    94, 1, 1, 1, 96, 288, 1, 97, 1, 96, 1, 1, 97, 96, 1, 96, 1, 48, 1, 96, 
    96, 1, 1, 96, 1, 1, 1, 48, 1, 43, 1, 1, 48, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 48, 1, 48, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 
    1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 48, 96, 1, 1, 96, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 48, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 48, 96, 48, 1, 
    288, 1, 288, 1, 96, 288, 1, 288, 1, 1, 288, 1, 93, 288, 1, 288, 1, 288, 
    1, 288, 1, 1, 288, 1, 288, 288, 1, 1, 288, 1, 288, 1, 96, 1, 96, 96, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 48, 1, 96, 1, 90, 
    96, 96, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 48, 1, 48, 1, 95, 96, 1, 96, 
    1, 1, 96, 1, 48, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 48, 1, 48, 1, 96, 96, 1, 48, 1, 1, 1, 96, 1, 1, 96, 1, 1, 95, 
    288, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 93, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 95, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 24, 96, 1, 1, 96, 1, 1, 22, 1, 96, 1, 24, 24, 1, 
    96, 1, 96, 1, 96, 96, 1, 24, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 94, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 49, 96, 1, 1, 1, 1, 96, 
    288, 48, 1, 1, 288, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    9, 96, 1, 288, 1, 288, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 24, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 288, 1, 96, 288, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 288, 1, 1, 1, 1, 96, 1, 1, 1, 288, 
    96, 1, 135, 1, 1, 1, 96, 1, 288, 1, 141, 96, 1, 1, 34, 1, 1, 1, 1, 95, 1, 
    1, 96, 288, 1, 1, 96, 1, 96, 1, 1, 1, 93, 1, 1, 1, 96, 288, 1, 288, 1, 1, 
    1, 288, 1, 1, 96, 1, 1, 288, 1, 1, 1, 1, 288, 1, 1, 288, 1, 1, 1, 24, 1, 
    1, 24, 1, 1, 1, 96, 288, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 288, 264, 1, 1, 287, 1, 1, 1, 1, 96, 96, 96, 1, 96, 1, 96, 
    288, 1, 96, 96, 1, 96, 273, 1, 96, 1, 96, 1, 1, 96, 24, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 24, 24, 96, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 48, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 92, 1, 96, 1, 96, 96, 
    96, 1, 96, 1, 96, 96, 1, 1, 120, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 105, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 
    1, 1, 92, 1, 96, 1, 1, 96, 240, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 96, 1, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 120, 240, 96, 1, 120, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 
    45, 1, 1, 1, 1, 240, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 288, 1, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 
    1, 48, 1, 24, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 95, 1, 48, 
    48, 1, 1, 1, 97, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 96, 1, 96, 1, 48, 1, 1, 96, 96, 1, 93, 1, 1, 1, 1, 48, 1, 
    48, 48, 1, 48, 1, 1, 48, 1, 96, 48, 1, 96, 1, 1, 96, 1, 48, 1, 96, 1, 96, 
    1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 48, 1, 96, 288, 1, 1, 96, 1, 48, 1, 96, 
    1, 96, 1, 96, 1, 288, 1, 96, 1, 96, 1, 288, 1, 1, 96, 1, 1, 48, 1, 288, 
    96, 1, 288, 144, 1, 96, 1, 1, 1, 48, 1, 48, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 99, 1, 99, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 48, 1, 96, 1, 97, 96, 1, 1, 96, 1, 96, 48, 1, 
    96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 94, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 98, 96, 96, 1, 
    96, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 288, 1, 288, 1, 1, 96, 1, 94, 1, 96, 96, 1, 96, 96, 1, 96, 1, 
    81, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 
    96, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 
    1, 96, 96, 96, 96, 1, 96, 96, 96, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 
    1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 96, 1, 96, 1, 26, 1, 96, 96, 96, 1, 
    96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 96, 96, 1, 
    96, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 96, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 18, 1, 96, 1, 96, 1, 95, 1, 1, 1, 96, 96, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 96, 96, 1, 96, 96, 96, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 
    96, 96, 96, 1, 96, 1, 89, 96, 1, 96, 96, 1, 1, 96, 92, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 
    1, 96, 48, 1, 48, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 96, 1, 96, 96, 96, 1, 96, 96, 1, 24, 96, 1, 96, 96, 1, 1, 
    96, 96, 1, 96, 1, 96, 1, 96, 1, 48, 1, 1, 96, 1, 48, 1, 96, 96, 1, 96, 1, 
    96, 1, 25, 1, 25, 96, 96, 1, 88, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 96, 1, 1, 47, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    96, 1, 96, 1, 1, 96, 96, 96, 1, 1, 96, 96, 96, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 82, 1, 96, 1, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 96, 96, 
    96, 1, 1, 1, 96, 92, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 14, 96, 1, 1, 1, 24, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 95, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 
    96, 96, 96, 96, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    288, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 88, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 
    1, 87, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 96, 96, 1, 144, 96, 1, 1, 144, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 288, 1, 96, 1, 96, 1, 1, 96, 1, 288, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 288, 96, 288, 1, 1, 96, 1, 1, 288, 1, 1, 96, 1, 1, 1, 288, 1, 
    1, 96, 1, 1, 1, 189, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 144, 1, 96, 1, 96, 1, 96, 1, 288, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 
    1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 90, 1, 96, 1, 96, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 95, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 96, 96, 1, 96, 1, 96, 1, 96, 1, 81, 1, 96, 1, 
    96, 1, 96, 96, 1, 82, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 96, 88, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 86, 96, 1, 1, 96, 37, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 94, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 90, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 92, 1, 96, 96, 
    1, 1, 1, 96, 8, 1, 1, 96, 1, 96, 1, 96, 1, 144, 1, 96, 1, 58, 96, 1, 1, 
    1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 48, 1, 96, 48, 
    1, 1, 1, 48, 96, 1, 47, 1, 1, 1, 46, 48, 1, 1, 48, 1, 48, 1, 48, 1, 48, 
    1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 96, 1, 48, 1, 288, 1, 1, 288, 1, 1, 96, 
    1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 95, 1, 95, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 95, 96, 288, 1, 1, 96, 
    96, 1, 96, 288, 1, 1, 96, 1, 288, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 288, 288, 288, 288, 
    288, 96, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1440, 1, 1, 1, 
    288, 96, 96, 1, 48, 1, 96, 96, 1, 1, 288, 1, 1, 1, 278, 96, 1, 96, 1, 1, 
    288, 1, 288, 1, 288, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 96, 96, 1, 96, 1, 288, 1, 96, 1, 1, 96, 96, 51, 95, 
    1, 1, 96, 1, 1, 96, 1, 96, 96, 96, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    24, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 96, 1, 1, 
    96, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 288, 1, 288, 1, 96, 1, 75, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 24, 24, 1, 190, 1, 1, 
    96, 1, 47, 48, 1, 48, 1, 96, 1, 286, 96, 1, 1, 96, 1, 1, 96, 93, 1, 96, 
    1, 96, 1, 94, 1, 1, 48, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 96, 1, 96, 95, 1, 96, 1, 96, 1, 1, 95, 1, 96, 1, 96, 1, 96, 
    46, 96, 1, 96, 48, 1, 96, 48, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 
    1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 93, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 69, 1, 49, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 
    76, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 95, 
    1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 62, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 34, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 35, 
    1, 1, 86, 1, 96, 96, 1, 1, 96, 1, 96, 1, 95, 1, 96, 88, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 94, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 50, 
    96, 1, 1, 96, 1, 96, 1, 73, 96, 1, 1, 57, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 95, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 
    37, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 95, 
    96, 1, 95, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 93, 1, 96, 1, 96, 1, 
    92, 1, 84, 1, 32, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 96, 1, 
    96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 288, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 288, 1, 1, 288, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 88, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 288, 1, 1, 
    1, 288, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 95, 1, 96, 
    1, 1, 96, 1, 1, 96, 96, 96, 94, 88, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 96, 96, 1, 96, 62, 62, 1, 96, 1, 1, 89, 1, 96, 1, 1, 96, 1, 1, 
    92, 1, 96, 1, 96, 96, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    87, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 95, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 14, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 289, 1, 96, 288, 96, 96, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 25, 1, 1, 96, 96, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 1, 84, 1, 
    96, 1, 96, 1, 38, 1, 91, 1, 99, 1, 96, 1, 81, 1, 95, 1, 33, 1, 1, 97, 1, 
    1, 94, 1, 91, 1, 93, 1, 1, 94, 1, 89, 1, 1, 88, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 88, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 288, 288, 1, 288, 
    1, 1, 96, 1, 1, 1, 288, 1, 288, 288, 1, 288, 1, 288, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 96, 1, 288, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 
    288, 1, 288, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 145, 1, 288, 267, 1, 96, 
    1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 1, 1, 29, 94, 1, 1, 96, 89, 1, 1, 96, 96, 1, 1, 95, 1, 96, 1, 96, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 95, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 96, 96, 1, 1, 96, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 90, 1, 96, 1, 71, 
    1, 1, 95, 1, 1, 96, 96, 96, 1, 96, 1, 96, 1, 52, 1, 1, 96, 96, 1, 96, 96, 
    1, 1, 96, 49, 1, 95, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 288, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 288, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    96, 96, 1, 96, 96, 1, 96, 80, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 94, 96, 1, 96, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 94, 96, 1, 1, 96, 1, 1, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 96, 1, 95, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 92, 96, 1, 
    96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 
    1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 96, 45, 96, 1, 1, 96, 81, 
    1, 96, 1, 1, 96, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 24, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 88, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 90, 288, 1, 288, 4, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 94, 1, 83, 96, 96, 1, 96, 1, 1, 1, 96, 89, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 92, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 69, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 54, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 36, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 1, 96, 1, 94, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 97, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 96, 1, 1, 94, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 288, 1, 288, 1, 1, 288, 1, 264, 1, 1, 
    1, 92, 288, 1, 1, 1, 96, 288, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 288, 288, 1, 288, 1, 1, 288, 1, 288, 1, 1, 1, 288, 1, 24, 
    1, 1, 1, 281, 1, 288, 1, 1, 288, 1, 287, 1, 288, 1, 288, 1, 288, 1, 1, 
    24, 1, 1, 288, 285, 1, 288, 1, 288, 264, 1, 288, 1, 288, 1, 288, 1, 1, 
    288, 288, 1, 288, 264, 1, 290, 1, 1, 288, 288, 1, 1, 288, 1, 1, 96, 48, 
    1, 1, 96, 1, 1, 1, 48, 1, 1, 96, 47, 1, 1, 48, 1, 96, 48, 1, 1, 1, 94, 
    48, 1, 1, 1, 264, 288, 1, 48, 1, 288, 1, 288, 1, 1, 288, 1, 288, 1, 1, 
    255, 287, 1, 48, 1, 96, 1, 46, 1, 1, 1, 1, 96, 96, 46, 1, 1, 1, 96, 94, 
    1, 1, 96, 1, 24, 24, 1, 96, 1, 96, 1, 46, 24, 1, 96, 96, 1, 96, 1, 96, 
    48, 1, 24, 24, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    1, 48, 24, 1, 96, 1, 61, 1, 96, 1, 48, 48, 1, 48, 1, 48, 1, 24, 1, 48, 1, 
    1, 1, 24, 1, 1, 96, 277, 1, 1, 1, 1, 89, 1, 24, 288, 1, 1, 288, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 288, 1, 96, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 22, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 95, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 98, 96, 1, 1, 47, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 92, 1, 1, 1, 1, 55, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 24, 96, 1, 1, 24, 24, 1, 
    286, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 
    156, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 96, 1, 96, 1, 1, 1, 85, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 86, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 96, 96, 96, 96, 1, 96, 1, 96, 96, 96, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 96, 1, 24, 1, 1, 1, 24, 1, 1, 
    1, 24, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 
    1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 96, 96, 1, 96, 1, 1, 96, 1, 48, 48, 1, 
    1, 96, 1, 48, 1, 1, 24, 1, 1, 1, 48, 96, 1, 1, 1, 48, 1, 96, 1, 96, 48, 
    1, 1, 48, 1, 1, 48, 1, 24, 1, 24, 1, 96, 1, 1, 1, 48, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 24, 1, 1, 48, 1, 1, 96, 1, 92, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 24, 24, 96, 1, 96, 1, 1, 96, 48, 1, 1, 96, 1, 
    48, 1, 1, 48, 1, 96, 1, 1, 48, 1, 1, 96, 1, 1, 26, 1, 1, 1, 1, 96, 1, 96, 
    1, 48, 1, 48, 1, 1, 1, 96, 84, 48, 1, 1, 24, 95, 1, 24, 1, 96, 96, 1, 1, 
    96, 96, 96, 1, 70, 1, 48, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    24, 1, 1, 96, 1, 24, 1, 1, 96, 1, 1, 48, 24, 1, 1, 96, 96, 1, 1, 92, 1, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 94, 1, 96, 1, 1, 24, 1, 1, 96, 1, 
    1, 48, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 23, 
    1, 96, 1, 48, 1, 1, 96, 1, 1, 94, 1, 1, 48, 1, 1, 96, 1, 1, 1, 1, 48, 1, 
    48, 1, 1, 96, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 96, 1, 96, 1, 96, 288, 
    1, 1, 96, 1, 1, 1, 1, 290, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 24, 1, 
    1, 1, 96, 96, 1, 1, 96, 1, 48, 1, 1, 96, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 
    48, 1, 96, 1, 1, 1, 48, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 92, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 288, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 48, 48, 1, 1, 48, 48, 1, 1, 24, 
    1, 288, 24, 1, 48, 1, 48, 1, 96, 1, 1, 1, 48, 1, 48, 1, 1, 96, 1, 1, 1, 
    48, 1, 1, 96, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 24, 1, 24, 1, 48, 1, 1, 
    48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 96, 24, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 48, 1, 1, 48, 1, 24, 1, 1, 48, 1, 1, 1, 48, 48, 1, 96, 
    1, 1, 48, 1, 1, 96, 96, 1, 48, 1, 48, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 24, 24, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 93, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 24, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    73, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 24, 24, 1, 24, 96, 1, 1, 1, 288, 1, 96, 1, 1, 96, 1, 96, 
    96, 24, 30, 1, 24, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 92, 1, 
    96, 96, 1, 24, 1, 96, 24, 1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 24, 27, 90, 15, 1, 1, 96, 1, 24, 24, 1, 1, 96, 24, 1, 96, 1, 96, 
    1, 96, 1, 24, 96, 1, 1, 1, 1, 96, 1, 1, 86, 1, 1, 60, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 62, 1, 96, 1, 1, 96, 1, 1, 96, 1, 48, 1, 1, 
    1, 48, 48, 1, 1, 24, 1, 1, 96, 1, 48, 1, 1, 48, 1, 1, 1, 48, 1, 48, 1, 1, 
    1, 96, 96, 1, 1, 1, 48, 1, 96, 1, 1, 48, 1, 48, 1, 1, 48, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 62, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 93, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 48, 
    1, 1, 1, 1, 37, 48, 1, 1, 96, 1, 1, 24, 1, 1, 96, 1, 1, 48, 1, 1, 1, 48, 
    1, 48, 1, 1, 96, 1, 1, 95, 1, 1, 96, 1, 1, 24, 1, 96, 1, 48, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 48, 96, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 24, 144, 1, 
    1, 1, 24, 1, 23, 96, 1, 1, 1, 24, 48, 1, 1, 48, 96, 1, 1, 48, 1, 24, 1, 
    96, 1, 1, 46, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 48, 1, 48, 1, 24, 1, 48, 
    1, 1, 24, 1, 1, 1, 1, 48, 96, 24, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 24, 1, 
    24, 1, 1, 48, 1, 1, 1, 1, 24, 1, 96, 1, 1, 96, 88, 48, 1, 1, 48, 1, 1, 
    48, 1, 1, 48, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 90, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 48, 1, 96, 96, 96, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 24, 48, 96, 96, 
    23, 24, 24, 1, 96, 1, 46, 48, 96, 96, 48, 24, 24, 24, 96, 1, 48, 96, 48, 
    288, 96, 96, 1, 96, 24, 1, 48, 48, 1, 48, 48, 48, 24, 1, 96, 96, 96, 1, 
    1, 1, 1, 96, 1, 1, 285, 288, 1, 1, 288, 1, 1, 96, 1, 96, 96, 1, 1, 288, 
    1, 1, 96, 1, 1, 1, 288, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 24, 1, 
    1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 95, 1, 96, 1, 
    1, 1, 96, 1, 24, 24, 1, 96, 1, 1, 1, 50, 1, 1, 1, 96, 1, 1, 48, 96, 1, 1, 
    1, 48, 48, 48, 24, 24, 1, 1, 24, 96, 1, 48, 48, 1, 96, 1, 48, 1, 1, 48, 
    48, 1, 48, 48, 1, 48, 24, 96, 1, 1, 1, 1, 96, 48, 48, 48, 1, 96, 1, 96, 
    1, 96, 96, 1, 1, 1, 24, 24, 96, 1, 1, 1, 48, 1, 1, 24, 1, 1, 48, 24, 1, 
    1, 240, 1, 1, 1, 1, 24, 1, 1, 96, 24, 96, 1, 96, 56, 1, 96, 1, 48, 1, 96, 
    1, 96, 1, 96, 1, 48, 1, 1, 1, 1, 96, 48, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 48, 1, 96, 1, 1, 96, 1, 48, 1, 1, 48, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 48, 1, 96, 1, 48, 1, 1, 48, 96, 48, 1, 48, 1, 1, 1, 1, 96, 1, 
    96, 1, 96, 96, 1, 96, 4, 1, 96, 96, 1, 96, 1, 96, 1, 96, 48, 1, 48, 1, 
    48, 96, 1, 1, 48, 1, 1, 96, 48, 1, 48, 1, 1, 1, 33, 1, 48, 48, 1, 48, 1, 
    48, 1, 48, 1, 96, 1, 96, 96, 1, 36, 1, 1, 1, 24, 1, 1, 24, 1, 1, 240, 1, 
    1, 1, 1, 96, 24, 1, 1, 24, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 96, 96, 96, 1, 
    1, 1, 1, 1, 240, 1, 1, 24, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 96, 1, 
    1, 1, 96, 1, 1, 56, 1, 24, 96, 48, 48, 1, 1, 96, 96, 48, 1, 96, 1, 96, 
    96, 240, 96, 1, 1, 48, 96, 1, 48, 48, 96, 1, 96, 96, 1, 96, 48, 1, 48, 
    96, 1, 1, 1, 1, 48, 1, 96, 240, 1, 1, 1, 1, 24, 1, 1, 1, 48, 1, 48, 1, 1, 
    1, 40, 1, 1, 48, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 96, 1, 48, 1, 1, 1, 
    24, 1, 1, 1, 1, 24, 1, 1, 24, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 95, 1, 1, 96, 96, 1, 85, 1, 1, 1, 96, 1, 48, 1, 96, 1, 
    1, 1, 1, 90, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 95, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 73, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 72, 1, 96, 
    96, 1, 94, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 94, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 95, 1, 96, 1, 
    96, 96, 1, 96, 96, 1, 1, 1, 1, 95, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 87, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 
    96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 96, 96, 1, 1, 60, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 90, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 95, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 95, 
    1, 1, 288, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 288, 1, 1, 1, 1, 95, 96, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 288, 1, 1, 1, 96, 1, 1, 1, 96, 1, 288, 288, 288, 
    1, 288, 288, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    95, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 288, 1, 1, 288, 1, 1, 95, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    288, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 
    1, 96, 1, 96, 96, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 
    1, 95, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 288, 1, 288, 1, 1, 1, 96, 1, 1, 
    288, 1, 1, 288, 1, 1, 96, 1, 96, 1, 288, 1, 1, 288, 1, 1, 96, 1, 288, 1, 
    288, 1, 288, 1, 288, 1, 288, 1, 288, 1, 288, 1, 288, 288, 1, 1, 96, 1, 1, 
    288, 1, 288, 1, 1, 288, 288, 1, 288, 1, 1, 288, 288, 1, 288, 1, 288, 1, 
    1, 1, 1, 1, 288, 1, 288, 1, 288, 1, 288, 1, 1, 196, 288, 1, 1, 288, 288, 
    1, 1, 288, 288, 1, 1, 288, 1, 288, 1, 288, 1, 288, 1, 288, 288, 1, 288, 
    96, 1, 1, 288, 1, 288, 1, 1, 288, 288, 1, 1, 96, 96, 1, 1, 96, 96, 96, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 93, 1, 96, 1, 1, 1, 96, 96, 96, 1, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 95, 1, 
    96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 68, 1, 1, 96, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    96, 96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 92, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 95, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 46, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 11, 96, 1, 
    1, 288, 1, 96, 1, 1, 96, 1, 1, 96, 1, 288, 1, 288, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 93, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 16, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 96, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 144, 1, 1, 1, 
    96, 1, 288, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 95, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 
    1, 1, 64, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 288, 288, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 80, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 93, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 93, 1, 96, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 288, 96, 1, 1, 96, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 94, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 94, 1, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 96, 1, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 90, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 91, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 96, 1, 96, 1, 94, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    101, 1, 101, 1, 93, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 94, 
    96, 1, 1, 1, 96, 1, 96, 1, 23, 1, 1, 96, 94, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 95, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 95, 1, 96, 96, 96, 
    1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 192, 96, 1, 192, 1, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 
    1, 96, 1, 94, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 95, 96, 1, 96, 1, 96, 1, 96, 96, 96, 96, 1, 
    96, 1, 96, 1, 81, 1, 96, 1, 44, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 96, 1, 1, 65, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 119, 1, 
    1, 96, 1, 95, 1, 1, 96, 1, 96, 1, 48, 98, 98, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 95, 1, 164, 1, 164, 1, 96, 1, 
    96, 1, 1, 94, 97, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 100, 1, 96, 1, 1, 96, 1, 99, 
    1, 96, 96, 1, 1, 96, 1, 1, 97, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 97, 1, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 24, 24, 1, 
    24, 96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 94, 83, 1, 96, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 62, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    94, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 92, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 92, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 
    1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 
    96, 1, 1, 96, 1, 96, 96, 1, 35, 1, 1, 43, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    96, 1, 96, 76, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    80, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 
    1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 24, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 95, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    89, 1, 96, 1, 76, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 85, 1, 96, 1, 96, 
    1, 96, 1, 62, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 90, 96, 1, 96, 94, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 
    1, 96, 1, 95, 1, 96, 91, 1, 95, 96, 96, 1, 96, 1, 96, 1, 100, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 98, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 94, 1, 96, 
    1, 288, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 288, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 93, 1, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 49, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 288, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 94, 1, 1, 95, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 85, 1, 85, 1, 85, 1, 85, 85, 1, 1, 86, 1, 1, 82, 1, 82, 82, 1, 
    1, 1, 1, 82, 1, 82, 1, 82, 1, 86, 1, 1, 1, 96, 1, 96, 96, 1, 1, 86, 1, 
    86, 1, 86, 1, 1, 87, 1, 59, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 93, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 84, 1, 1, 1, 84, 1, 84, 1, 78, 96, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 35, 1, 40, 96, 1, 96, 1, 96, 1, 
    1, 1, 84, 1, 84, 1, 1, 84, 1, 1, 84, 1, 1, 1, 84, 1, 1, 1, 96, 1, 96, 96, 
    1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 84, 96, 1, 89, 1, 96, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 1, 42, 1, 1, 96, 1, 96, 1, 96, 96, 96, 1, 96, 96, 1, 1, 1, 
    96, 1, 96, 96, 1, 1, 96, 96, 96, 1, 1, 96, 20, 1, 1, 96, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 144, 1, 1, 1, 48, 1, 
    96, 1, 1, 96, 1, 1, 96, 227, 1, 1, 1, 48, 96, 96, 1, 1, 96, 1, 1, 1, 1, 
    144, 1, 144, 1, 144, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 91, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 53, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 96, 96, 1, 48, 1, 96, 1, 96, 1, 1, 96, 1, 48, 1, 96, 96, 1, 96, 1, 
    96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 1, 96, 1, 96, 96, 
    1, 96, 1, 96, 96, 1, 96, 49, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 32, 1, 86, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 96, 96, 96, 48, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 24, 1, 96, 1, 24, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 24, 1, 48, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 96, 96, 1, 96, 96, 96, 1, 96, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 95, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 
    94, 1, 96, 1, 66, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 93, 1, 96, 96, 1, 96, 1, 96, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 
    96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 56, 1, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 288, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 96, 1, 
    96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 97, 1, 96, 1, 1, 95, 1, 96, 96, 1, 96, 96, 97, 97, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 72, 1, 96, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 81, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 89, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 97, 1, 
    96, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 96, 96, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 56, 84, 1, 1, 96, 1, 96, 96, 1, 
    1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 96, 1, 96, 1, 1, 
    1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 99, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 41, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 52, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    96, 1, 28, 28, 1, 96, 1, 96, 1, 1, 96, 1, 44, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 1, 86, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 48, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 
    1, 96, 1, 96, 96, 96, 1, 89, 1, 48, 1, 1, 1, 1, 48, 96, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 112, 1, 1, 96, 96, 1, 1, 1, 96, 1, 108, 1, 104, 1, 1, 98, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 95, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 67, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 96, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 97, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 1, 114, 1, 
    1, 108, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 106, 1, 96, 1, 1, 1, 96, 
    1, 1, 112, 1, 96, 1, 1, 107, 1, 131, 1, 101, 1, 127, 1, 137, 1, 1, 126, 
    1, 128, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 96, 96, 1, 1, 96, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 1, 
    96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 94, 1, 1, 1, 96, 1, 96, 1, 1, 97, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 96, 
    96, 1, 96, 1, 1, 288, 97, 1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    95, 1, 1, 96, 1, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 96, 96, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    1, 96, 1, 96, 96, 96, 96, 1, 1, 48, 1, 96, 1, 1, 42, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 87, 1, 96, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 96, 96, 1, 1, 1, 88, 
    1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 51, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 24, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 64, 
    1, 64, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 96, 1, 96, 1, 96, 96, 1, 96, 
    1, 96, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    96, 1, 1, 94, 1, 96, 1, 96, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 113, 1, 96, 96, 1, 96, 1, 96, 96, 1, 225, 1, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 112, 1, 96, 1, 102, 1, 100, 1, 96, 1, 96, 1, 288, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 52, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 96, 96, 96, 1, 1, 96, 91, 1, 1, 96, 1, 1, 1, 96, 96, 96, 96, 
    96, 96, 1, 1, 24, 24, 96, 96, 96, 96, 96, 96, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 96, 96, 96, 96, 96, 
    96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 1, 96, 1, 96, 96, 
    1, 96, 1, 96, 96, 96, 96, 96, 96, 96, 95, 96, 96, 96, 96, 96, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 
    1, 1, 24, 1, 1, 48, 48, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 48, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 48, 1, 48, 
    1, 24, 1, 1, 35, 1, 1, 186, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 24, 1, 96, 1, 1, 1, 1, 96, 48, 1, 1, 96, 96, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    91, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 84, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 58, 1, 48, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 137, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 88, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 71, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 288, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 96, 
    96, 1, 96, 1, 1, 1, 24, 24, 1, 1440, 1, 24, 24, 1, 24, 24, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 890, 1, 1, 96, 1, 1, 96, 
    1, 89, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 288, 1, 1211, 
    1, 1, 96, 1, 1, 1, 1, 96, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 88, 1, 96, 1, 96, 
    1, 1, 1, 1, 288, 288, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    95, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1 ;

 v00010_validated =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 144, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 87, 1, 1, 1, 
    97, 1, 95, 1, 1, 1, 1, 1, 144, 1, 1, 1, 111, 1, 1, 1, 144, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 26, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 144, 
    1, 1, 1, 1, 144, 1, 1, 144, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 
    1, 1, 96, 1, 1, 144, 1, 1, 1, 1, 144, 1, 1, 144, 1, 1, 1, 1, 1, 144, 1, 
    144, 1, 1, 1, 1, 144, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 93, 1, 1, 1, 1, 1, 93, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 240, 1, 226, 1, 1, 1, 1, 
    1, 240, 1, 240, 1, 1, 1, 240, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 120, 1, 
    240, 1, 1, 1, 240, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 52, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 24, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 24, 1, 1, 1, 1, 1, 20, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 1, 
    24, 1, 1, 1, 24, 1, 1, 120, 1, 1, 1, 1, 1, 24, 23, 1, 1, 120, 1, 1, 1, 1, 
    120, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 24, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 24, 1, 20, 1, 24, 1, 24, 1, 24, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 
    48, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 27, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 47, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 25, 1, 1, 1, 48, 1, 1, 1, 1, 
    48, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 46, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 231, 1, 1, 240, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 208, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 48, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 96, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 
    1, 288, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 92, 92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 103, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 24, 24, 1, 1, 1, 24, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 96, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 13, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    84, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 95, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 93, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 95, 1, 1, 1, 1, 61, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 93, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 73, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 84, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 93, 1, 1, 95, 1, 1, 61, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    91, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 96, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 89, 1, 1, 1, 1, 96, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 95, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 94, 1, 95, 1, 1, 95, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 61, 1, 61, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 82, 1, 1, 1, 1, 1, 94, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 91, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 32, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 93, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 14, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 90, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 84, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 36, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 92, 1, 1, 1, 
    94, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 95, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 48, 1, 1, 1, 24, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 24, 1, 1, 1, 1, 96, 1, 1, 24, 1, 24, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 24, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 24, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 70, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 91, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 288, 1, 1, 
    1, 289, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 34, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 
    289, 1, 1, 1, 1, 1, 1, 192, 1, 1, 1, 288, 1, 1, 1, 288, 1, 1, 1, 288, 1, 
    1, 24, 1, 1, 1, 24, 1, 1, 1, 288, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 24, 1, 1, 24, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    24, 1, 1, 24, 1, 1, 24, 24, 24, 24, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 276, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 120, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 289, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 46, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 76, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 3, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 78, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    86, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 288, 1, 1, 1, 1, 
    288, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 144, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 288, 1, 1, 1, 96, 1, 1, 1, 288, 1, 1, 96, 1, 1, 189, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 25, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 89, 1, 1, 1, 1, 1, 95, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1440, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    97, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 51, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 35, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 36, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 21, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 47, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    22, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 92, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    22, 1, 1, 11, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 276, 276, 276, 276, 276, 276, 276, 276, 1, 1, 
    276, 276, 276, 276, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 72, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 50, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 48, 1, 1, 23, 1, 1, 48, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 24, 1, 1, 25, 1, 1, 1, 
    1, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 24, 1, 1, 1, 1, 
    1, 24, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 48, 96, 1, 1, 96, 1, 1, 96, 1, 72, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    94, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 93, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 45, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 67, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 25, 1, 25, 1, 25, 1, 25, 1, 
    1, 1, 1, 1, 1, 1, 144, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 42, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 5, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 18, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 95, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 93, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 85, 1, 20, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 94, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 82, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 90, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 24, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 96, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 84, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    84, 1, 1, 1, 1, 1, 83, 1, 1, 1, 1, 1, 84, 1, 1, 1, 84, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 95, 1, 1, 1, 1, 144, 1, 1, 1, 1, 1, 1, 1, 96, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 24, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 78, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 73, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 96, 
    1, 1, 1, 1, 1, 1, 98, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 86, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 97, 1, 1, 1, 1, 1, 1, 1, 1, 96, 114, 
    1, 1, 108, 1, 1, 1, 1, 96, 1, 1, 1, 1, 87, 1, 1, 106, 1, 1, 1, 1, 96, 96, 
    1, 1, 96, 1, 1, 113, 1, 107, 1, 1, 1, 1, 101, 1, 1, 1, 1, 1, 126, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 25, 
    1, 1, 1, 1, 1, 24, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 49, 1, 
    1, 1, 48, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 96, 1, 97, 1, 1, 96, 1, 1, 96, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 96, 1, 1, 1, 48, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 40, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 24, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 64, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 47, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    96, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 91, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 96, 96, 96, 96, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 25, 25, 25, 25, 25, 25, 25, 
    25, 25, 25, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 93, 1, 93, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 95, 1, 95, 1, 95, 24, 1, 24, 1, 1, 24, 1, 24, 1, 1, 1, 24, 
    1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 24, 1, 1, 24, 1, 1, 
    1, 48, 24, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 48, 1, 24, 1, 1, 96, 1, 24, 1, 
    24, 1, 24, 1, 24, 1, 1, 24, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 48, 1, 48, 1, 24, 1, 
    1, 60, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 48, 1, 48, 1, 96, 1, 1, 24, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 24, 1, 24, 94, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    49, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 96, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 18, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 
    48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 85, 85, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 88, 
    1, 1, 85, 1, 1, 23, 1, 19, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 24, 1, 
    24, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 92, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    720, 720, 720, 720, 720, 720, 720, 720, 720, 720, 720, 720, 720, 720, 
    720, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 24, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 24, 24, 1, 1, 24, 1, 1, 1, 24, 
    1, 1, 1, 24, 1, 24, 1, 24, 1, 95, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 96, 1, 1, 90, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 82, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 52, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 35, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 19, 1, 19, 19, 23, 21, 24, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    24, 1, 24, 1, 1, 24, 1, 24, 6, 1, 8, 1, 19, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 10, 10, 1, 1, 23, 1, 5, 1, 18, 18, 1, 19, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1 ;

 v00095_validated =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 144, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 78, 1, 97, 1, 
    1, 1, 95, 1, 1, 1, 1, 1, 144, 1, 1, 1, 96, 1, 1, 1, 144, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    37, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 144, 1, 
    1, 1, 1, 144, 1, 1, 144, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 144, 1, 1, 96, 
    1, 1, 1, 1, 144, 1, 1, 1, 1, 144, 1, 1, 144, 1, 1, 1, 144, 1, 1, 1, 144, 
    1, 1, 144, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    93, 1, 1, 1, 1, 1, 93, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 240, 1, 226, 1, 1, 1, 1, 1, 240, 1, 
    240, 1, 1, 1, 240, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 120, 1, 240, 1, 1, 1, 
    240, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 24, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 27, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 46, 1, 1, 1, 1, 1, 47, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 25, 1, 1, 1, 48, 1, 1, 48, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 231, 1, 1, 240, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 205, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 288, 1, 1, 
    1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 92, 92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 48, 1, 1, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 84, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 95, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 92, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 58, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    93, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 73, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 84, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 
    1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 90, 1, 1, 1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 89, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 88, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 94, 1, 95, 1, 1, 1, 1, 95, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 60, 1, 61, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 86, 1, 1, 1, 1, 94, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 91, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 32, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    93, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 84, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 12, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 22, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 36, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 92, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 90, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 
    289, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 289, 1, 1, 
    1, 1, 1, 1, 192, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 288, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 276, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 120, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 289, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 46, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 84, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 
    1, 288, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 44, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 67, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 97, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 83, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 21, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 22, 1, 1, 11, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 88, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 44, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 
    1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    73, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 50, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 23, 1, 1, 48, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 24, 1, 1, 25, 1, 1, 1, 1, 1, 
    24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 24, 1, 1, 1, 24, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 
    1, 24, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    1, 1, 96, 48, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 93, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 44, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 69, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 25, 1, 25, 1, 25, 1, 25, 1, 1, 1, 
    1, 1, 1, 1, 144, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 5, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 18, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 85, 1, 13, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    82, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 90, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 84, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 84, 1, 1, 1, 1, 1, 83, 1, 1, 1, 1, 1, 84, 1, 1, 1, 84, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 41, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 25, 1, 1, 
    1, 1, 1, 24, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 49, 1, 1, 1, 
    48, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 50, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 52, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 96, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    91, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 93, 1, 92, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 95, 1, 95, 1, 95, 1, 1, 24, 1, 24, 24, 1, 1, 1, 24, 1, 1, 1, 
    24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 1, 24, 1, 24, 1, 1, 24, 1, 
    1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 96, 1, 24, 
    1, 24, 1, 24, 1, 24, 1, 1, 24, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    60, 1, 1, 1, 1, 1, 24, 1, 1, 96, 48, 1, 48, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 24, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 96, 31, 1, 1, 1, 
    1, 24, 24, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 18, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    96, 1, 1, 85, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 88, 85, 1, 1, 23, 1, 19, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 24, 1, 24, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 92, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 24, 1, 1, 1, 24, 1, 24, 1, 24, 1, 95, 1, 24, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 88, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    82, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 24, 1, 24, 1, 1, 1, 1, 1, 6, 1, 8, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1 ;

 v00035_validated =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 90, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 36, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 15, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 276, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 33, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 12, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 65, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 22, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 48, 48, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 56, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 48, 
    1, 1, 1, 1, 1, 1, 45, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 48, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 24, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 7, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 25, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    19, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 v00036_validated =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 240, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 90, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 34, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 15, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 276, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 36, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    65, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 25, 25, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 52, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 44, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 24, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 716, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 24, 
    1, 24, 24, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 7, 1, 1, 1, 1, 1, 1, 1, 1, 1, 25, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 19, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 v00045_validated =
  96, 45, 96, 96, 1, 96, 96, 24, 24, 96, 48, 48, 96, 96, 96, 96, 96, 96, 96, 
    96, 24, 96, 96, 96, 48, 96, 24, 144, 96, 48, 96, 96, 96, 96, 48, 24, 96, 
    96, 96, 96, 96, 96, 96, 96, 96, 96, 142, 96, 96, 96, 144, 96, 24, 96, 96, 
    96, 144, 96, 24, 96, 144, 96, 144, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 95, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 43, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    240, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 90, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 288, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 288, 
    1, 1, 1, 1, 96, 288, 1, 1, 96, 1, 1, 1, 288, 1, 1, 1, 96, 96, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 95, 1, 1, 1, 1, 69, 1, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 95, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 93, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 94, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 85, 1, 1, 1, 85, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 95, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 92, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 86, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 42, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 92, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 48, 1, 1, 48, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 96, 48, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 48, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 89, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 288, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 93, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 42, 1, 1, 
    96, 1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 24, 1, 96, 1, 1, 1, 288, 1, 1, 96, 1, 96, 1, 
    1, 96, 1, 96, 1, 1, 1, 288, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 
    288, 1, 1, 264, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 288, 1, 1, 288, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 288, 
    1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 288, 1, 1, 93, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 
    1, 24, 1, 1, 1, 96, 1, 1, 24, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 288, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 92, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 48, 1, 1, 1, 48, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 
    48, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 
    1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 48, 1, 288, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 48, 1, 288, 1, 1, 1, 1, 1, 1, 1, 
    1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 48, 1, 1, 1, 43, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 48, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 288, 1, 1, 288, 1, 1, 288, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 288, 1, 288, 1, 1, 288, 1, 288, 288, 1, 96, 1, 1, 288, 1, 288, 1, 
    288, 1, 288, 288, 1, 288, 1, 1, 288, 288, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 288, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 24, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 135, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 7, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 
    95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 288, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 288, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 43, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 288, 1, 
    1, 288, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 95, 1, 96, 1, 1, 1, 1, 1, 
    1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 68, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 89, 
    1, 1, 1, 77, 1, 91, 1, 96, 1, 1, 1, 89, 1, 92, 1, 1, 62, 1, 1, 95, 1, 93, 
    1, 93, 1, 1, 92, 1, 92, 1, 1, 93, 1, 1, 4, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 56, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 48, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 47, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 22, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 40, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 92, 1, 1, 1, 1, 54, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 279, 1, 1, 
    1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 288, 1, 1, 288, 1, 1, 1, 1, 1, 
    1, 288, 1, 1, 288, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 
    1, 1, 24, 1, 1, 1, 96, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 48, 1, 96, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 96, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 92, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 48, 1, 1, 
    96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 96, 1, 1, 96, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    96, 1, 1, 48, 1, 1, 48, 1, 1, 24, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 48, 1, 1, 96, 1, 1, 24, 1, 1, 96, 1, 48, 1, 1, 1, 48, 1, 48, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 
    1, 48, 1, 1, 1, 1, 96, 1, 96, 1, 1, 48, 1, 1, 96, 1, 1, 48, 1, 1, 48, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 96, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 24, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 96, 1, 88, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 24, 1, 1, 1, 96, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 92, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    24, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 44, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 48, 48, 1, 1, 1, 48, 1, 1, 24, 1, 
    1, 1, 1, 48, 1, 1, 48, 48, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 96, 1, 
    1, 1, 24, 24, 1, 1, 96, 1, 1, 1, 1, 1, 24, 1, 96, 1, 24, 1, 1, 96, 1, 1, 
    96, 1, 24, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 24, 1, 1, 96, 1, 
    24, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 
    1, 1, 96, 1, 1, 24, 1, 1, 96, 1, 1, 48, 48, 1, 1, 1, 1, 48, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 24, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 1, 1, 144, 1, 1, 23, 1, 1, 1, 1, 24, 1, 
    1, 1, 48, 1, 1, 1, 144, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 
    1, 96, 1, 1, 1, 48, 1, 1, 1, 1, 1, 24, 1, 1, 48, 1, 24, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 24, 1, 1, 48, 1, 1, 48, 1, 1, 48, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 50, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 55, 1, 96, 1, 48, 1, 1, 1, 96, 1, 
    96, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 48, 1, 
    1, 1, 96, 96, 1, 96, 1, 96, 1, 1, 48, 1, 96, 1, 96, 1, 96, 1, 96, 1, 48, 
    1, 96, 1, 1, 48, 1, 1, 1, 48, 1, 48, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 71, 1, 1, 96, 1, 96, 1, 96, 1, 1, 48, 1, 48, 1, 1, 1, 96, 1, 48, 96, 
    1, 1, 48, 1, 48, 1, 1, 1, 33, 1, 1, 48, 1, 48, 1, 48, 1, 48, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 
    1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 56, 1, 96, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 88, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 
    96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 95, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 
    1, 1, 1, 1, 1, 95, 1, 1, 1, 96, 1, 96, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 48, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 96, 1, 95, 1, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 96, 1, 
    1, 96, 288, 1, 1, 288, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 96, 1, 1, 1, 1, 288, 1, 1, 1, 96, 1, 1, 288, 1, 1, 288, 1, 1, 96, 
    1, 1, 1, 288, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1378, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 
    288, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 
    1, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 48, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 
    1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 29, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 31, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 48, 1, 1, 96, 1, 1, 92, 1, 
    1, 96, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 288, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 
    1, 80, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 94, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 118, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 98, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    96, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 92, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 
    1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 44, 1, 1, 
    1, 48, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 
    1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 48, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 48, 1, 
    1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 
    48, 1, 48, 1, 48, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 48, 
    1, 1, 1, 48, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 32, 1, 1, 48, 1, 1, 48, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 91, 288, 96, 96, 
    96, 96, 96, 96, 1, 96, 96, 1, 1, 96, 96, 96, 96, 96, 96, 1, 96, 96, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 
    96, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 96, 1, 1, 1, 1, 274, 96, 96, 96, 
    1, 1, 96, 1, 1, 96, 96, 96, 96, 1, 1, 96, 1, 1, 96, 96, 1, 1, 1, 96, 1, 
    96, 48, 1, 1, 96, 1, 1, 1, 96, 98, 288, 17, 288, 96, 96, 1, 96, 96, 96, 
    99, 96, 96, 96, 96, 96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 
    1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 96, 96, 1, 1, 24, 96, 96, 1, 96, 1, 96, 
    96, 126, 126, 1, 96, 126, 96, 96, 96, 72, 96, 96, 48, 96, 263, 1, 1, 1, 
    1, 1, 1, 264, 96, 96, 96, 96, 96, 96, 96, 288, 96, 288, 288, 288, 288, 
    288, 288, 288, 288, 288, 288, 288, 288, 288, 288, 288, 96, 96, 288, 288, 
    288, 288, 288, 288, 288, 288, 288, 288, 288, 288, 1, 1, 288, 288, 288, 
    288, 288, 48, 288, 288, 288, 288, 288, 288, 288, 288, 48, 288, 288, 288, 
    288, 288, 288, 288, 288, 288, 288, 288, 288, 288, 1, 1, 288, 288, 288, 
    288, 288, 288, 288, 288, 1, 1, 288, 288, 288, 288, 288, 288, 288, 96, 48, 
    288, 1, 96, 288, 288, 288, 96, 96, 1, 1, 288, 288, 288, 1, 1, 288, 288, 
    288, 1, 288, 288, 288, 288, 96, 288, 288, 288, 288, 288, 288, 288, 96, 1, 
    1, 1, 1, 96, 96, 1, 1, 288, 96, 1, 96, 96, 48, 288, 288, 1, 1, 1, 288, 1, 
    1, 96, 96, 96, 38, 96, 1, 96, 48, 96, 48, 1, 1, 96, 48, 48, 1, 48, 96, 1, 
    1, 48, 48, 48, 96, 48, 96, 48, 96, 48, 288, 96, 48, 96, 288, 48, 1, 1, 1, 
    288, 288, 1, 1, 1, 1, 1, 288, 1, 1, 48, 48, 96, 1, 1, 1, 1, 1, 1, 48, 1, 
    1, 1, 1, 1, 1, 1, 96, 48, 96, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 96, 
    96, 48, 1, 96, 1, 1, 48, 288, 1, 1, 1, 1, 288, 48, 1, 1, 1, 1, 48, 96, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 48, 48, 1, 1, 48, 288, 96, 
    96, 1, 1, 288, 1, 1, 1, 288, 288, 288, 149, 96, 96, 1, 1, 48, 96, 96, 96, 
    24, 288, 1, 1, 1, 1, 48, 24, 288, 96, 96, 48, 96, 96, 1, 1, 288, 48, 1, 
    1, 96, 48, 48, 96, 48, 96, 1, 1, 96, 96, 48, 1, 1, 1, 1, 96, 24, 96, 1, 
    1, 48, 1, 96, 1, 288, 288, 288, 288, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 24, 48, 1, 1, 96, 1, 1, 96, 1, 1, 1, 96, 48, 96, 1, 24, 288, 1, 1, 96, 
    48, 1, 1, 288, 1, 1, 1, 1, 48, 96, 288, 288, 96, 1, 1, 288, 1, 1, 1, 1, 
    89, 96, 95, 1, 1, 1, 1, 1, 288, 1, 1, 96, 96, 96, 96, 1, 1, 48, 96, 96, 
    288, 1, 1, 24, 1, 1, 96, 1, 1, 1, 288, 1, 1, 48, 96, 96, 96, 48, 96, 96, 
    96, 96, 96, 1, 1, 96, 1, 1, 96, 96, 96, 96, 96, 96, 1, 96, 96, 96, 96, 
    96, 96, 96, 1, 1, 1, 1, 96, 1, 96, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 96, 1, 96, 96, 1, 96, 1, 1, 96, 96, 
    96, 96, 1, 1, 96, 96, 1, 1, 1, 96, 96, 1, 96, 96, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 96, 96, 96, 96, 96, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 2, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 
    96, 96, 1, 1, 1, 144, 96, 1, 1, 24, 288, 1, 1, 288, 1, 1, 48, 96, 1, 96, 
    96, 24, 48, 96, 96, 1, 96, 1, 1, 48, 1, 1, 1, 96, 96, 96, 48, 96, 96, 1, 
    1, 1, 1, 48, 1, 1, 48, 96, 55, 1, 1, 288, 288, 1, 288, 288, 96, 288, 149, 
    96, 1, 1, 48, 288, 288, 288, 288, 48, 48, 1, 1, 273, 288, 288, 288, 48, 
    288, 1, 1, 48, 288, 1, 1, 288, 96, 1, 1, 288, 48, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 96, 1, 1, 1, 1, 96, 96, 96, 1, 288, 1, 1, 1, 1, 1, 96, 1, 1, 
    96, 96, 232, 1, 1, 1, 1, 96, 288, 1, 1, 45, 1, 1, 96, 96, 1, 1, 1, 1, 96, 
    1, 24, 96, 96, 1, 1, 24, 1, 96, 1, 1, 24, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 
    96, 96, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 890, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 96, 96, 1, 1, 96, 1, 1, 1, 1, 1440, 1, 1, 96, 
    24, 96, 1, 1, 1, 1, 96, 96, 1, 78, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 96, 1, 
    1, 1, 24, 1, 1, 96, 1, 1, 1, 96, 1, 1, 96, 96, 96, 96, 96, 96, 96, 96, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 80, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 144, 144, 144, 144, 96, 144, 
    144, 144, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 10, 11, 1, 23, 1, 4, 
    1, 1, 18, 1, 18, 144, 144, 96, 1, 96, 144, 1, 1, 96 ;

 v00062_validated =
  1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 91, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 20, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 48, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 86, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 48, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 288, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 24, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 23, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 96, 96, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 56, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 96, 1, 1, 96, 1, 1, 96, 1, 1, 
    96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    92, 1, 1, 1, 1, 24, 1, 96, 96, 96, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 96, 
    96, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 96, 1, 1, 1, 96, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 96, 96, 1, 1, 96, 96, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1378, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 71, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 95, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 112, 1, 1, 1, 1, 1, 1, 1, 1, 1, 108, 1, 104, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 131, 1, 1, 1, 127, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 91, 
    1, 1, 1, 1, 1, 1, 1, 1, 76, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 92, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 
    96, 1, 96, 1, 96, 1, 96, 1, 1, 96, 96, 1, 96, 1, 96, 1, 96, 1, 96, 1, 96, 
    1, 96, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 v00054_validated =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 95, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 23, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 1, 48, 1, 1, 
    1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 48, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 48, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 56, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 71, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 46, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 96, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 24, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 96, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 96, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 24, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 v00060_description =
  "USGS:02339495:00011:00002",
  "USGS:02339495:00011:00001",
  "USGS:02342500:00011:00001",
  "USGS:02342500:00011:00002",
  "USGS:0234296910:00011:00002",
  "USGS:023432415:00011:00016",
  "USGS:023432415:00011:00003",
  "USGS:023432415:00011:00002",
  "USGS:023432415:00011:00001",
  "USGS:023432415:00011:00017",
  "USGS:023432415:00011:00018",
  "USGS:02361000:00011:00010",
  "USGS:02361000:00011:00011",
  "USGS:02361000:00011:00002",
  "USGS:02361000:00011:00003",
  "USGS:02361500:00011:00005",
  "USGS:02361500:00011:00006",
  "USGS:02361500:00011:00001",
  "USGS:02361500:00011:00002",
  "USGS:02362000:00011:00002",
  "USGS:02362240:00011:00001",
  "USGS:02362240:00011:00002",
  "USGS:02363000:00011:00001",
  "USGS:02363000:00011:00002",
  "USGS:02364000:00011:00001",
  "USGS:02364500:00011:00005",
  "USGS:02364500:00011:00006",
  "USGS:02364500:00011:00001",
  "USGS:02364500:00011:00002",
  "USGS:02369800:00011:00002",
  "USGS:02369800:00011:00003",
  "USGS:02371500:00011:00005",
  "USGS:02371500:00011:00006",
  "USGS:02372250:00011:00001",
  "USGS:02372250:00011:00002",
  "USGS:02372422:00011:00005",
  "USGS:02372422:00011:00004",
  "USGS:02372430:00011:00003",
  "USGS:02372430:00011:00001",
  "USGS:02373000:00011:00001",
  "USGS:02373000:00011:00002",
  "USGS:02374250:00011:00002",
  "USGS:02374250:00011:00001",
  "USGS:02374500:00011:00001",
  "USGS:02374500:00011:00002",
  "USGS:02374700:00011:00004",
  "USGS:02374700:00011:00002",
  "USGS:02374700:00011:00001",
  "USGS:02374745:00011:00002",
  "USGS:02374745:00011:00001",
  "USGS:02374950:00011:00002",
  "USGS:02374950:00011:00001",
  "USGS:02376500:00011:00002",
  "USGS:02376500:00011:00001",
  "USGS:02377560:00011:00001",
  "USGS:02377570:00011:00002",
  "USGS:02377570:00011:00001",
  "USGS:02377750:00011:00001",
  "USGS:02378170:00011:00002",
  "USGS:02378170:00011:00001",
  "USGS:02378300:00011:00002",
  "USGS:02378300:00011:00001",
  "USGS:02378500:00011:00003",
  "USGS:02378500:00011:00001",
  "USGS:02378500:00011:00002",
  "USGS:02397530:00011:00001",
  "USGS:02397530:00011:00007",
  "USGS:02397530:00011:00026",
  "USGS:02397530:00011:00027",
  "USGS:02397530:00011:00017",
  "USGS:02397530:00011:00002",
  "USGS:02397530:00011:00003",
  "USGS:02397530:00011:00004",
  "USGS:02398300:00011:00001",
  "USGS:02398300:00011:00002",
  "USGS:02399200:00011:00001",
  "USGS:02399200:00011:00002",
  "USGS:02399500:00011:00002",
  "USGS:02400100:00011:00001",
  "USGS:02400100:00011:00002",
  "USGS:02400496:00011:00002",
  "USGS:02400500:00011:00003",
  "USGS:02400680:00011:00002",
  "USGS:02400680:00011:00001",
  "USGS:02401000:00011:00001",
  "USGS:02401000:00011:00002",
  "USGS:02401390:00011:00001",
  "USGS:02401390:00011:00002",
  "USGS:02401895:00011:00002",
  "USGS:02401895:00011:00001",
  "USGS:02403310:00011:00001",
  "USGS:07176321:00011:00002",
  "USGS:02404400:00011:00001",
  "USGS:02404400:00011:00002",
  "USGS:02405500:00011:00004",
  "USGS:02405500:00011:00001",
  "USGS:02405500:00011:00002",
  "USGS:02406500:00011:00001",
  "USGS:02406500:00011:00002",
  "USGS:02406930:00011:00002",
  "USGS:02406930:00011:00001",
  "USGS:02407000:00011:00004",
  "USGS:02407000:00011:00002",
  "USGS:02407000:00011:00003",
  "USGS:02407514:00011:00004",
  "USGS:02407514:00011:00002",
  "USGS:02407514:00011:00001",
  "USGS:02407526:00011:00001",
  "USGS:02408150:00011:00001",
  "USGS:02408540:00011:00001",
  "USGS:02408540:00011:00002",
  "USGS:01118300:00011:00004",
  "USGS:01118300:00011:00016",
  "USGS:01118300:00011:00001",
  "USGS:01118300:00011:00003",
  "USGS:01119382:00011:00013",
  "USGS:01119382:00011:00015",
  "USGS:01119382:00011:00009",
  "USGS:01119382:00011:00002",
  "USGS:01119382:00011:00001",
  "USGS:01119500:00011:00002",
  "USGS:01119500:00011:00005",
  "USGS:01120790:00011:00004",
  "USGS:01120790:00011:00005",
  "USGS:01120790:00011:00007",
  "USGS:01120790:00011:00001",
  "USGS:01120790:00011:00002",
  "USGS:01121000:00011:00001",
  "USGS:01121000:00011:00003",
  "USGS:01121330:00011:00001",
  "USGS:01121330:00011:00002",
  "USGS:01121500:00011:00002",
  "USGS:02471078:00011:00002",
  "USGS:02471078:00011:00001",
  "USGS:02479945:00011:00002",
  "USGS:02479945:00011:00001",
  "USGS:02479980:00011:00002",
  "USGS:02479980:00011:00001",
  "USGS:02480002:00011:00002",
  "USGS:02480002:00011:00001",
  "USGS:03572690:00011:00002",
  "USGS:03572690:00011:00001",
  "USGS:03574500:00011:00004",
  "USGS:03574500:00011:00005",
  "USGS:0357479650:00011:00001",
  "USGS:03575100:00011:00002",
  "USGS:03575100:00011:00001",
  "USGS:0357526200:00011:00003",
  "USGS:0357526200:00011:00002",
  "USGS:0357526200:00011:00001",
  "USGS:03575272:00011:00004",
  "USGS:03575272:00011:00002",
  "USGS:03575272:00011:00001",
  "USGS:03575500:00011:00002",
  "USGS:0357568650:00011:00003",
  "USGS:0357568650:00011:00002",
  "USGS:0357568650:00011:00001",
  "USGS:0357568980:00011:00003",
  "USGS:0357568980:00011:00002",
  "USGS:0357568980:00011:00001",
  "USGS:03575700:00011:00001",
  "USGS:03575700:00011:00002",
  "USGS:03575700:00011:00003",
  "USGS:03575830:00011:00001",
  "USGS:03575830:00011:00002",
  "USGS:03575830:00011:00003",
  "USGS:0357586650:00011:00003",
  "USGS:0357586650:00011:00002",
  "USGS:0357586650:00011:00001",
  "USGS:0357587090:00011:00003",
  "USGS:0357587090:00011:00002",
  "USGS:0357587090:00011:00001",
  "USGS:0357587140:00011:00003",
  "USGS:0357587140:00011:00002",
  "USGS:0357587140:00011:00001",
  "USGS:0357587400:00011:00003",
  "USGS:0357587400:00011:00002",
  "USGS:0357587400:00011:00001",
  "USGS:0357587728:00011:00001",
  "USGS:0357587728:00011:00002",
  "USGS:0357587728:00011:00003",
  "USGS:02411600:00011:00003",
  "USGS:03575890:00011:00001",
  "USGS:03575890:00011:00002",
  "USGS:03575890:00011:00003",
  "USGS:0357591500:00011:00003",
  "USGS:0357591500:00011:00002",
  "USGS:0357591500:00011:00001",
  "USGS:03575950:00011:00001",
  "USGS:03575950:00011:00002",
  "USGS:03575950:00011:00003",
  "USGS:03575980:00011:00001",
  "USGS:03575980:00011:00003",
  "USGS:03575980:00011:00002",
  "USGS:03576250:00011:00001",
  "USGS:03576250:00011:00002",
  "USGS:03576500:00011:00002",
  "USGS:03576500:00011:00003",
  "USGS:03577150:00011:00002",
  "USGS:03577225:00011:00002",
  "USGS:03577225:00011:00001",
  "USGS:03586500:00011:00002",
  "USGS:03586500:00011:00003",
  "USGS:03589500:00011:00003",
  "USGS:03590000:00011:00002",
  "USGS:03592500:00011:00003",
  "USGS:322047086214301:00011:00001",
  "USGS:322500085551201:00011:00001",
  "USGS:332934086353801:00011:00001",
  "USGS:333103086524501:00011:00001",
  "USGS:333204087324601:00011:00001",
  "USGS:333205086493701:00011:00002",
  "USGS:333437086430801:00011:00001",
  "USGS:335929087021001:00011:00001",
  "USGS:340618086344001:00011:00001",
  "USGS:342718087285601:00011:00001",
  "USGS:343843085403201:00011:00001",
  "USGS:02204520:00011:00015",
  "USGS:02204520:00011:00005",
  "USGS:02204520:00011:00016",
  "USGS:02204520:00011:00017",
  "USGS:02204520:00011:00002",
  "USGS:02204520:00011:00001",
  "USGS:02205000:00011:00006",
  "USGS:02205865:00011:00004",
  "USGS:02205865:00011:00003",
  "USGS:02205865:00011:00002",
  "USGS:02205865:00011:00001",
  "USGS:02205865:00011:00005",
  "USGS:02207120:00011:00006",
  "USGS:02207120:00011:00003",
  "USGS:02207120:00011:00002",
  "USGS:02207120:00011:00001",
  "USGS:02207120:00011:00007",
  "USGS:02207130:00011:00005",
  "USGS:02207130:00011:00004",
  "USGS:02207135:00011:00007",
  "USGS:02207135:00011:00005",
  "USGS:02207135:00011:00004",
  "USGS:02207135:00011:00008",
  "USGS:02207135:00011:00009",
  "USGS:02412000:00011:00001",
  "USGS:02412000:00011:00002",
  "USGS:02413300:00011:00001",
  "USGS:02413300:00011:00002",
  "USGS:02414500:00011:00001",
  "USGS:02414500:00011:00002",
  "USGS:02414715:00011:00001",
  "USGS:02414715:00011:00002",
  "USGS:02415000:00011:00001",
  "USGS:02415000:00011:00002",
  "USGS:02418230:00011:00002",
  "USGS:02418230:00011:00001",
  "USGS:02418760:00011:00002",
  "USGS:02418760:00011:00001",
  "USGS:02419000:00011:00001",
  "USGS:02419000:00011:00002",
  "USGS:02419500:00011:00002",
  "USGS:02419890:00011:00004",
  "USGS:02419890:00011:00002",
  "USGS:02419890:00011:00001",
  "USGS:02419890:00011:00006",
  "USGS:02419890:00011:00008",
  "USGS:02419988:00011:00001",
  "USGS:02420000:00011:00007",
  "USGS:02420000:00011:00003",
  "USGS:02420000:00011:00004",
  "USGS:02420490:00011:00001",
  "USGS:02421000:00011:00001",
  "USGS:02421000:00011:00002",
  "USGS:02421350:00011:00002",
  "USGS:02421350:00011:00001",
  "USGS:02421351:00011:00002",
  "USGS:02422500:00011:00001",
  "USGS:02422500:00011:00002",
  "USGS:02423000:00011:00003",
  "USGS:02423110:00011:00001",
  "USGS:02423110:00011:00003",
  "USGS:02423130:00011:00003",
  "USGS:02423130:00011:00002",
  "USGS:02423130:00011:00001",
  "USGS:02423130:00011:00004",
  "USGS:02423130:00011:00005",
  "USGS:02423160:00011:00003",
  "USGS:02423160:00011:00002",
  "USGS:02423160:00011:00001",
  "USGS:02423160:00011:00004",
  "USGS:02423160:00011:00005",
  "USGS:02423380:00011:00006",
  "USGS:02423380:00011:00007",
  "USGS:02423397:00011:00004",
  "USGS:02423397:00011:00002",
  "USGS:02423397:00011:00001",
  "USGS:02423397:00011:00005",
  "USGS:02423397:00011:00006",
  "USGS:02423400:00011:00004",
  "USGS:02423400:00011:00002",
  "USGS:02423414:00011:00002",
  "USGS:02423414:00011:00001",
  "USGS:02423425:00011:00002",
  "USGS:02423425:00011:00001",
  "USGS:07176321:00011:00001",
  "USGS:02423496:00011:00003",
  "USGS:02423496:00011:00002",
  "USGS:02423496:00011:00001",
  "USGS:02423496:00011:00004",
  "USGS:02423496:00011:00005",
  "USGS:02423500:00011:00001",
  "USGS:02423500:00011:00002",
  "USGS:0242354750:00011:00002",
  "USGS:0242354750:00011:00001",
  "USGS:02423555:00011:00002",
  "USGS:02423555:00011:00001",
  "USGS:02423630:00011:00001",
  "USGS:02423630:00011:00002",
  "USGS:02424000:00011:00004",
  "USGS:02424000:00011:00005",
  "USGS:02424590:00011:00001",
  "USGS:02425000:00011:00001",
  "USGS:02425000:00011:00002",
  "USGS:02427250:00011:00002",
  "USGS:02427250:00011:00001",
  "USGS:02427505:00011:00002",
  "USGS:02427505:00011:00001",
  "USGS:02427506:00011:00002",
  "USGS:02427830:00011:00002",
  "USGS:02427830:00011:00001",
  "USGS:02428400:00011:00002",
  "USGS:02428400:00011:00003",
  "USGS:02428400:00011:00006",
  "USGS:02428400:00011:00007",
  "USGS:02428400:00011:00008",
  "USGS:02428400:00011:00009",
  "USGS:02428400:00011:00010",
  "USGS:02428400:00011:00011",
  "USGS:02428401:00011:00002",
  "USGS:02438000:00011:00001",
  "USGS:02438000:00011:00002",
  "USGS:02444160:00011:00001",
  "USGS:02444160:00011:00003",
  "USGS:02444160:00011:00005",
  "USGS:02444160:00011:00006",
  "USGS:02444160:00011:00007",
  "USGS:02444160:00011:00008",
  "USGS:02444161:00011:00001",
  "USGS:02446500:00011:00001",
  "USGS:02446500:00011:00002",
  "USGS:02447025:00011:00001",
  "USGS:02447025:00011:00003",
  "USGS:02447025:00011:00005",
  "USGS:02447025:00011:00006",
  "USGS:02447025:00011:00007",
  "USGS:02447025:00011:00008",
  "USGS:02447025:00011:00009",
  "USGS:02447026:00011:00001",
  "USGS:02448500:00011:00001",
  "USGS:02448500:00011:00002",
  "USGS:02448900:00011:00002",
  "USGS:02448900:00011:00001",
  "USGS:02449882:00011:00002",
  "USGS:02449882:00011:00001",
  "USGS:02193340:00011:00001",
  "USGS:02193340:00011:00002",
  "USGS:15085100:00011:00007",
  "USGS:15085100:00011:00002",
  "USGS:15085100:00011:00005",
  "USGS:15099900:00011:00013",
  "USGS:15099900:00011:00015",
  "USGS:15099900:00011:00001",
  "USGS:15099900:00011:00002",
  "USGS:15099900:00011:00003",
  "USGS:15100000:00011:00012",
  "USGS:15100000:00011:00001",
  "USGS:15100000:00011:00002",
  "USGS:15100000:00011:00003",
  "USGS:15101490:00011:00002",
  "USGS:15101490:00011:00003",
  "USGS:15129120:00011:00005",
  "USGS:15129120:00011:00015",
  "USGS:15129120:00011:00016",
  "USGS:15129120:00011:00003",
  "USGS:15129120:00011:00001",
  "USGS:15129120:00011:00002",
  "USGS:15129120:00011:00006",
  "USGS:15129500:00011:00008",
  "USGS:15129500:00011:00002",
  "USGS:15129500:00011:00019",
  "USGS:15129500:00011:00004",
  "USGS:15129500:00011:00006",
  "USGS:15129500:00011:00009",
  "USGS:15200280:00011:00001",
  "USGS:15200280:00011:00002",
  "USGS:15200280:00011:00003",
  "USGS:15214000:00011:00016",
  "USGS:15214000:00011:00017",
  "USGS:15214000:00011:00020",
  "USGS:15214000:00011:00005",
  "USGS:15214000:00011:00002",
  "USGS:15214000:00011:00003",
  "USGS:15225997:00011:00001",
  "USGS:15225997:00011:00002",
  "USGS:15225997:00011:00005",
  "USGS:15226620:00011:00002",
  "USGS:15226620:00011:00001",
  "USGS:15236895:00011:00002",
  "USGS:15236895:00011:00004",
  "USGS:15236895:00011:00025",
  "USGS:15236895:00011:00014",
  "USGS:15236895:00011:00016",
  "USGS:15236895:00011:00020",
  "USGS:15236895:00011:00026",
  "USGS:15236895:00011:00019",
  "USGS:15236895:00011:00001",
  "USGS:15236895:00011:00023",
  "USGS:15236900:00011:00005",
  "USGS:15236900:00011:00016",
  "USGS:15236900:00011:00001",
  "USGS:15236900:00011:00003",
  "USGS:15237730:00011:00003",
  "USGS:15237730:00011:00014",
  "USGS:15237730:00011:00001",
  "USGS:15238648:00011:00003",
  "USGS:15238648:00011:00004",
  "USGS:15238648:00011:00001",
  "USGS:15238648:00011:00002",
  "USGS:15238648:00011:00008",
  "USGS:15238990:00011:00004",
  "USGS:15238990:00011:00002",
  "USGS:15238990:00011:00007",
  "USGS:15238990:00011:00009",
  "USGS:15239001:00011:00004",
  "USGS:15239001:00011:00020",
  "USGS:15239001:00011:00021",
  "USGS:15239001:00011:00019",
  "USGS:15239001:00011:00005",
  "USGS:15239001:00011:00018",
  "USGS:15239001:00011:00002",
  "USGS:15239001:00011:00001",
  "USGS:15239001:00011:00017",
  "USGS:15239001:00011:00007",
  "USGS:15239050:00011:00005",
  "USGS:15239050:00011:00001",
  "USGS:15239050:00011:00002",
  "USGS:15239050:00011:00008",
  "USGS:15239060:00011:00004",
  "USGS:15239060:00011:00002",
  "USGS:15239060:00011:00001",
  "USGS:15239060:00011:00007",
  "USGS:15239070:00011:00002",
  "USGS:15239070:00011:00007",
  "USGS:15239070:00011:00003",
  "USGS:15239070:00011:00005",
  "USGS:15239070:00011:00014",
  "USGS:15239070:00011:00006",
  "USGS:15239900:00011:00004",
  "USGS:15239900:00011:00002",
  "USGS:15243900:00011:00005",
  "USGS:15243900:00011:00001",
  "USGS:15243900:00011:00003",
  "USGS:15258000:00011:00003",
  "USGS:15258000:00011:00017",
  "USGS:15258000:00011:00006",
  "USGS:15258000:00011:00004",
  "USGS:15258000:00011:00002",
  "USGS:15261000:00011:00003",
  "USGS:15261000:00011:00001",
  "USGS:15261000:00011:00002",
  "USGS:15266110:00011:00003",
  "USGS:15266110:00011:00002",
  "USGS:15266110:00011:00001",
  "USGS:15266300:00011:00017",
  "USGS:15266300:00011:00023",
  "USGS:15266300:00011:00001",
  "USGS:15266300:00011:00005",
  "USGS:15271000:00011:00015",
  "USGS:15271000:00011:00004",
  "USGS:15271000:00011:00005",
  "USGS:15274600:00011:00006",
  "USGS:15274600:00011:00005",
  "USGS:15275100:00011:00010",
  "USGS:15275100:00011:00007",
  "USGS:15276000:00011:00008",
  "USGS:15276000:00011:00002",
  "USGS:15276000:00011:00004",
  "USGS:15278000:00011:00002",
  "USGS:15278000:00011:00001",
  "USGS:15283700:00011:00014",
  "USGS:15283700:00011:00001",
  "USGS:15283700:00011:00002",
  "USGS:15284000:00011:00001",
  "USGS:15284000:00011:00002",
  "USGS:15284000:00011:00006",
  "USGS:15290000:00011:00003",
  "USGS:15290000:00011:00014",
  "USGS:15291700:00011:00012",
  "USGS:15291700:00011:00017",
  "USGS:15291700:00011:00001",
  "USGS:15291700:00011:00002",
  "USGS:15292000:00011:00005",
  "USGS:15292000:00011:00020",
  "USGS:15292000:00011:00001",
  "USGS:15292400:00011:00001",
  "USGS:15292400:00011:00002",
  "USGS:15292400:00011:00003",
  "USGS:15292400:00011:00013",
  "USGS:15292700:00011:00001",
  "USGS:15292700:00011:00019",
  "USGS:15292700:00011:00008",
  "USGS:15292700:00011:00002",
  "USGS:15292700:00011:00003",
  "USGS:15292700:00011:00020",
  "USGS:15292780:00011:00004",
  "USGS:15292780:00011:00005",
  "USGS:15292780:00011:00006",
  "USGS:15292780:00011:00015",
  "USGS:15292780:00011:00003",
  "USGS:15292800:00011:00016",
  "USGS:15292800:00011:00003",
  "USGS:15292800:00011:00006",
  "USGS:15292800:00011:00001",
  "USGS:15293200:00011:00013",
  "USGS:15293200:00011:00014",
  "USGS:15293200:00011:00003",
  "USGS:15293200:00011:00001",
  "USGS:15293200:00011:00002",
  "USGS:15293700:00011:00003",
  "USGS:15293700:00011:00001",
  "USGS:15293700:00011:00002",
  "USGS:15294005:00011:00017",
  "USGS:15294005:00011:00003",
  "USGS:15294005:00011:00006",
  "USGS:15294005:00011:00002",
  "USGS:15295700:00011:00004",
  "USGS:15295700:00011:00022",
  "USGS:15295700:00011:00018",
  "USGS:15295700:00011:00015",
  "USGS:15295700:00011:00016",
  "USGS:15297610:00011:00003",
  "USGS:15297610:00011:00001",
  "USGS:15297610:00011:00002",
  "USGS:15298040:00011:00001",
  "USGS:15298040:00011:00019",
  "USGS:15298040:00011:00002",
  "USGS:15298040:00011:00003",
  "USGS:15298040:00011:00017",
  "USGS:15300100:00011:00003",
  "USGS:15300100:00011:00013",
  "USGS:15300100:00011:00001",
  "USGS:15300100:00011:00002",
  "USGS:15300250:00011:00014",
  "USGS:15300250:00011:00016",
  "USGS:15300250:00011:00003",
  "USGS:15300250:00011:00001",
  "USGS:15300250:00011:00013",
  "USGS:15300300:00011:00014",
  "USGS:15300300:00011:00016",
  "USGS:15300300:00011:00012",
  "USGS:15300300:00011:00002",
  "USGS:15300300:00011:00013",
  "USGS:15302000:00011:00016",
  "USGS:15302000:00011:00018",
  "USGS:15302000:00011:00014",
  "USGS:15302000:00011:00004",
  "USGS:15302000:00011:00005",
  "USGS:01096000:00011:00001",
  "USGS:01096000:00011:00003",
  "USGS:01122000:00011:00001",
  "USGS:01122000:00011:00005",
  "USGS:01122500:00011:00001",
  "USGS:01122500:00011:00003",
  "USGS:01123000:00011:00001",
  "USGS:01123000:00011:00003",
  "USGS:011230695:00011:00002",
  "USGS:011230695:00011:00014",
  "USGS:01124000:00011:00001",
  "USGS:01124000:00011:00003",
  "USGS:01124151:00011:00014",
  "USGS:01124151:00011:00013",
  "USGS:01124151:00011:00001",
  "USGS:01124151:00011:00005",
  "USGS:01125100:00011:00002",
  "USGS:01125100:00011:00001",
  "USGS:01125490:00011:00001",
  "USGS:01125490:00011:00002",
  "USGS:01125500:00011:00004",
  "USGS:01125500:00011:00005",
  "USGS:01127000:00011:00002",
  "USGS:01127000:00011:00005",
  "USGS:01127500:00011:00016",
  "USGS:01127500:00011:00001",
  "USGS:01127500:00011:00006",
  "USGS:011277905:00011:00002",
  "USGS:011277905:00011:00001",
  "USGS:01184000:00011:00002",
  "USGS:01184000:00011:00005",
  "USGS:01184100:00011:00017",
  "USGS:01184100:00011:00019",
  "USGS:01184100:00011:00001",
  "USGS:01184100:00011:00007",
  "USGS:01184490:00011:00001",
  "USGS:01184490:00011:00004",
  "USGS:01186000:00011:00002",
  "USGS:01186000:00011:00005",
  "USGS:01186500:00011:00001",
  "USGS:01186500:00011:00004",
  "USGS:01187300:00011:00005",
  "USGS:01187300:00011:00006",
  "USGS:01187300:00011:00001",
  "USGS:01187300:00011:00002",
  "USGS:01188000:00011:00002",
  "USGS:01188000:00011:00004",
  "USGS:01188090:00011:00002",
  "USGS:01188090:00011:00003",
  "USGS:01189213:00011:00001",
  "USGS:01189995:00011:00002",
  "USGS:01189995:00011:00005",
  "USGS:01190070:00011:00005",
  "USGS:01191000:00011:00001",
  "USGS:01191000:00011:00002",
  "USGS:01192500:00011:00002",
  "USGS:01192500:00011:00014",
  "USGS:01192883:00011:00016",
  "USGS:01192883:00011:00018",
  "USGS:01192883:00011:00001",
  "USGS:01192883:00011:00006",
  "USGS:01193050:00011:00006",
  "USGS:01193050:00011:00026",
  "USGS:01193050:00011:00035",
  "USGS:01193050:00011:00012",
  "USGS:01193050:00011:00011",
  "USGS:01193050:00011:00009",
  "USGS:01193050:00011:00007",
  "USGS:01193050:00011:00010",
  "USGS:01193050:00011:00038",
  "USGS:01193050:00011:00037",
  "USGS:01193050:00011:00041",
  "USGS:01193500:00011:00001",
  "USGS:01193500:00011:00011",
  "USGS:01193500:00011:00002",
  "USGS:01193500:00011:00003",
  "USGS:01194000:00011:00005",
  "USGS:01194000:00011:00004",
  "USGS:01194000:00011:00001",
  "USGS:01194000:00011:00002",
  "USGS:01194500:00011:00017",
  "USGS:01194500:00011:00016",
  "USGS:01194500:00011:00003",
  "USGS:01194500:00011:00001",
  "USGS:01194500:00011:00002",
  "USGS:01194750:00011:00003",
  "USGS:01194750:00011:00010",
  "USGS:01194750:00011:00013",
  "USGS:01194750:00011:00001",
  "USGS:01194750:00011:00004",
  "USGS:01194750:00011:00011",
  "USGS:01194750:00011:00014",
  "USGS:01194750:00011:00006",
  "USGS:01194750:00011:00007",
  "USGS:01194750:00011:00008",
  "USGS:01194750:00011:00009",
  "USGS:01194750:00011:00005",
  "USGS:01194750:00011:00012",
  "USGS:01194750:00011:00015",
  "USGS:01194796:00011:00004",
  "USGS:01194796:00011:00006",
  "USGS:01194796:00011:00001",
  "USGS:01194796:00011:00005",
  "USGS:01194796:00011:00007",
  "USGS:01194796:00011:00009",
  "USGS:01194796:00011:00010",
  "USGS:01195100:00011:00004",
  "USGS:01195100:00011:00001",
  "USGS:01195100:00011:00003",
  "USGS:01195490:00011:00011",
  "USGS:01195490:00011:00002",
  "USGS:01195490:00011:00003",
  "USGS:01196500:00011:00001",
  "USGS:01196500:00011:00017",
  "USGS:01196500:00011:00014",
  "USGS:01196500:00011:00002",
  "USGS:01196500:00011:00003",
  "USGS:01196500:00011:00004",
  "USGS:01196500:00011:00016",
  "USGS:01196561:00011:00002",
  "USGS:01196561:00011:00001",
  "USGS:01196620:00011:00001",
  "USGS:01196620:00011:00003",
  "USGS:01199000:00011:00019",
  "USGS:01199000:00011:00018",
  "USGS:01199000:00011:00002",
  "USGS:01199000:00011:00003",
  "USGS:01199050:00011:00001",
  "USGS:01199050:00011:00003",
  "USGS:01200500:00011:00002",
  "USGS:01200500:00011:00008",
  "USGS:02457595:00011:00005",
  "USGS:01200600:00011:00002",
  "USGS:01200600:00011:00009",
  "USGS:01200600:00011:00003",
  "USGS:01200600:00011:00011",
  "USGS:01201487:00011:00014",
  "USGS:01201487:00011:00017",
  "USGS:01201487:00011:00003",
  "USGS:01201487:00011:00002",
  "USGS:01201487:00011:00001",
  "USGS:01201487:00011:00015",
  "USGS:01201487:00011:00016",
  "USGS:01202501:00011:00014",
  "USGS:01202501:00011:00002",
  "USGS:01202501:00011:00001",
  "USGS:012035055:00011:00002",
  "USGS:012035055:00011:00001",
  "USGS:01203510:00011:00001",
  "USGS:01203510:00011:00002",
  "USGS:01203600:00011:00001",
  "USGS:01203600:00011:00003",
  "USGS:01203805:00011:00019",
  "USGS:01203805:00011:00018",
  "USGS:01203805:00011:00001",
  "USGS:01203805:00011:00003",
  "USGS:01204000:00011:00002",
  "USGS:01204000:00011:00005",
  "USGS:07294800:00011:00001",
  "USGS:02450000:00011:00002",
  "USGS:02450000:00011:00003",
  "USGS:02450180:00011:00002",
  "USGS:02450180:00011:00003",
  "USGS:02450250:00011:00006",
  "USGS:02450250:00011:00001",
  "USGS:02450250:00011:00002",
  "USGS:02450825:00011:00002",
  "USGS:02450825:00011:00003",
  "USGS:02453000:00011:00003",
  "USGS:02453000:00011:00004",
  "USGS:02453500:00011:00009",
  "USGS:02453500:00011:00001",
  "USGS:02453500:00011:00002",
  "USGS:02454055:00011:00002",
  "USGS:02454055:00011:00001",
  "USGS:02455000:00011:00002",
  "USGS:02455000:00011:00003",
  "USGS:02455185:00011:00002",
  "USGS:02455185:00011:00001",
  "USGS:02455980:00011:00003",
  "USGS:02455980:00011:00001",
  "USGS:02455980:00011:00002",
  "USGS:02455980:00011:00004",
  "USGS:02455980:00011:00005",
  "USGS:02456500:00011:00002",
  "USGS:02456500:00011:00003",
  "USGS:02457000:00011:00002",
  "USGS:02457000:00011:00003",
  "USGS:02457595:00011:00003",
  "USGS:02457595:00011:00002",
  "USGS:02457595:00011:00001",
  "USGS:02457595:00011:00004",
  "USGS:02458148:00011:00004",
  "USGS:02458148:00011:00002",
  "USGS:02458148:00011:00001",
  "USGS:02458148:00011:00005",
  "USGS:02458190:00011:00002",
  "USGS:02458190:00011:00001",
  "USGS:02458300:00011:00003",
  "USGS:02458300:00011:00002",
  "USGS:02458450:00011:00004",
  "USGS:02458450:00011:00002",
  "USGS:02458450:00011:00003",
  "USGS:02458450:00011:00005",
  "USGS:02458450:00011:00006",
  "USGS:02458502:00011:00004",
  "USGS:02458502:00011:00002",
  "USGS:02458502:00011:00001",
  "USGS:02458502:00011:00005",
  "USGS:02458600:00011:00002",
  "USGS:02458600:00011:00001",
  "USGS:02461500:00011:00002",
  "USGS:02461500:00011:00003",
  "USGS:02462000:00011:00002",
  "USGS:02462000:00011:00003",
  "USGS:02462500:00011:00008",
  "USGS:02462500:00011:00003",
  "USGS:02462501:00011:00001",
  "USGS:02462951:00011:00005",
  "USGS:02462951:00011:00004",
  "USGS:02462952:00011:00001",
  "USGS:02464000:00011:00002",
  "USGS:02464000:00011:00003",
  "USGS:02464146:00011:00002",
  "USGS:02464146:00011:00001",
  "USGS:02464360:00011:00002",
  "USGS:02464360:00011:00003",
  "USGS:02464660:00011:00002",
  "USGS:02464660:00011:00001",
  "USGS:02464800:00011:00011",
  "USGS:02464800:00011:00003",
  "USGS:02464800:00011:00007",
  "USGS:02465000:00011:00003",
  "USGS:02465000:00011:00004",
  "USGS:02465005:00011:00001",
  "USGS:02465292:00011:00002",
  "USGS:02465292:00011:00001",
  "USGS:02465493:00011:00001",
  "USGS:02465493:00011:00002",
  "USGS:02466030:00011:00001",
  "USGS:02466030:00011:00003",
  "USGS:02466030:00011:00005",
  "USGS:02466030:00011:00006",
  "USGS:02466030:00011:00007",
  "USGS:02466030:00011:00008",
  "USGS:02466030:00011:00009",
  "USGS:02466030:00011:00010",
  "USGS:02466031:00011:00003",
  "USGS:02467000:00011:00001",
  "USGS:02467000:00011:00002",
  "USGS:02467001:00011:00002",
  "USGS:02467500:00011:00001",
  "USGS:02467500:00011:00002",
  "USGS:02469525:00011:00004",
  "USGS:02469525:00011:00001",
  "USGS:02469761:00011:00001",
  "USGS:02469761:00011:00002",
  "USGS:02469761:00011:00005",
  "USGS:02469761:00011:00006",
  "USGS:02469761:00011:00007",
  "USGS:02469761:00011:00008",
  "USGS:02469761:00011:00009",
  "USGS:02469761:00011:00010",
  "USGS:02469761:00011:00011",
  "USGS:02469761:00011:00012",
  "USGS:02469762:00011:00002",
  "USGS:02469800:00011:00001",
  "USGS:02469800:00011:00002",
  "USGS:02470050:00011:00001",
  "USGS:02470072:00011:00003",
  "USGS:02470072:00011:00002",
  "USGS:02470629:00011:00005",
  "USGS:02470629:00011:00004",
  "USGS:02470629:00011:00003",
  "USGS:02470629:00011:00026",
  "USGS:02470630:00011:00001",
  "USGS:02471001:00011:00001",
  "USGS:02471001:00011:00002",
  "USGS:02471019:00011:00002",
  "USGS:02471019:00011:00004",
  "USGS:03613000:00011:00003",
  "USGS:03613000:00011:00001",
  "USGS:01205500:00011:00002",
  "USGS:01205500:00011:00005",
  "USGS:01206900:00011:00001",
  "USGS:01206900:00011:00006",
  "USGS:01208011:00011:00002",
  "USGS:01208500:00011:00002",
  "USGS:01208500:00011:00003",
  "USGS:01208873:00011:00001",
  "USGS:01208873:00011:00002",
  "USGS:01208925:00011:00001",
  "USGS:01208925:00011:00002",
  "USGS:01208950:00011:00005",
  "USGS:01208950:00011:00006",
  "USGS:01208950:00011:00001",
  "USGS:01208950:00011:00003",
  "USGS:01208990:00011:00001",
  "USGS:01208990:00011:00003",
  "USGS:01209005:00011:00002",
  "USGS:01209005:00011:00001",
  "USGS:01209105:00011:00002",
  "USGS:01209105:00011:00001",
  "USGS:01209500:00011:00002",
  "USGS:01209500:00011:00003",
  "USGS:01209510:00011:00001",
  "USGS:012095493:00011:00001",
  "USGS:012095493:00011:00002",
  "USGS:01209700:00011:00001",
  "USGS:01209700:00011:00002",
  "USGS:01209761:00011:00002",
  "USGS:01209761:00011:00001",
  "USGS:01209788:00011:00001",
  "USGS:01209788:00011:00002",
  "USGS:01209901:00011:00001",
  "USGS:01209901:00011:00002",
  "USGS:01212500:00011:00003",
  "USGS:01212500:00011:00002",
  "USGS:01212500:00011:00001",
  "USGS:02176930:00011:00013",
  "USGS:02176930:00011:00003",
  "USGS:02176930:00011:00002",
  "USGS:02176930:00011:00001",
  "USGS:02178400:00011:00006",
  "USGS:02178400:00011:00002",
  "USGS:02178400:00011:00003",
  "USGS:02181350:00011:00005",
  "USGS:02181350:00011:00004",
  "USGS:02181350:00011:00001",
  "USGS:02181580:00011:00003",
  "USGS:02181580:00011:00002",
  "USGS:02181580:00011:00001",
  "USGS:02188600:00011:00005",
  "USGS:02188600:00011:00002",
  "USGS:02188600:00011:00003",
  "USGS:02191227:00011:00004",
  "USGS:02191227:00011:00001",
  "USGS:02191300:00011:00015",
  "USGS:02191300:00011:00013",
  "USGS:02191300:00011:00003",
  "USGS:15051010:00011:00003",
  "USGS:02191740:00011:00003",
  "USGS:02191740:00011:00002",
  "USGS:02191740:00011:00001",
  "USGS:02191743:00011:00003",
  "USGS:02191743:00011:00002",
  "USGS:02191743:00011:00001",
  "USGS:02192000:00011:00001",
  "USGS:02192000:00011:00002",
  "USGS:15008000:00011:00001",
  "USGS:15008000:00011:00002",
  "USGS:15009000:00011:00003",
  "USGS:15009000:00011:00014",
  "USGS:15009000:00011:00001",
  "USGS:15009000:00011:00002",
  "USGS:15009000:00011:00004",
  "USGS:15019990:00011:00002",
  "USGS:15019990:00011:00004",
  "USGS:15024800:00011:00019",
  "USGS:15024800:00011:00004",
  "USGS:15024800:00011:00002",
  "USGS:15024800:00011:00008",
  "USGS:15041200:00011:00016",
  "USGS:15041200:00011:00018",
  "USGS:15041200:00011:00020",
  "USGS:15041200:00011:00021",
  "USGS:15041200:00011:00017",
  "USGS:15041200:00011:00002",
  "USGS:15041200:00011:00005",
  "USGS:15041200:00011:00007",
  "USGS:15051010:00011:00014",
  "USGS:15051010:00011:00002",
  "USGS:15051010:00011:00005",
  "USGS:15052000:00011:00001",
  "USGS:15052000:00011:00002",
  "USGS:15052500:00011:00014",
  "USGS:15052500:00011:00003",
  "USGS:15052500:00011:00004",
  "USGS:15052500:00011:00005",
  "USGS:15055500:00011:00002",
  "USGS:15055500:00011:00001",
  "USGS:15056210:00011:00001",
  "USGS:15056210:00011:00002",
  "USGS:15056210:00011:00005",
  "USGS:15056210:00011:00003",
  "USGS:15056210:00011:00004",
  "USGS:15056500:00011:00008",
  "USGS:15056500:00011:00002",
  "USGS:15056500:00011:00006",
  "USGS:15056500:00011:00009",
  "USGS:15058700:00011:00001",
  "USGS:15058700:00011:00002",
  "USGS:15058700:00011:00003",
  "USGS:15072000:00011:00004",
  "USGS:15072000:00011:00001",
  "USGS:15072000:00011:00002",
  "USGS:15081497:00011:00006",
  "USGS:15081497:00011:00002",
  "USGS:15081497:00011:00004",
  "USGS:15081497:00011:00008",
  "USGS:410628073413301:00011:00001",
  "USGS:4121480721223:00011:00002",
  "USGS:4121480721223:00011:00003",
  "USGS:4121480721223:00011:00001",
  "USGS:412429073165101:00011:00002",
  "USGS:412825072410501:00011:00001",
  "USGS:412916073121701:00011:00001",
  "USGS:413535072253701:00011:00001",
  "USGS:414741072134501:00011:00001",
  "USGS:414831072173002:00011:00001",
  "USGS:02193500:00011:00014",
  "USGS:02193500:00011:00001",
  "USGS:02193500:00011:00004",
  "USGS:02195320:00011:00006",
  "USGS:02195320:00011:00004",
  "USGS:02195320:00011:00003",
  "USGS:02195520:00011:00001",
  "USGS:021964832:00011:00003",
  "USGS:021964832:00011:00005",
  "USGS:021964832:00011:00001",
  "USGS:02196485:00011:00004",
  "USGS:02196485:00011:00001",
  "USGS:02196835:00011:00003",
  "USGS:02196835:00011:00002",
  "USGS:02196835:00011:00001",
  "USGS:02196838:00011:00007",
  "USGS:02196838:00011:00006",
  "USGS:02196838:00011:00003",
  "USGS:02196838:00011:00004",
  "USGS:02196838:00011:00002",
  "USGS:02196838:00011:00018",
  "USGS:02196838:00011:00001",
  "USGS:02196999:00011:00002",
  "USGS:02196999:00011:00001",
  "USGS:02197000:00011:00001",
  "USGS:02197000:00011:00002",
  "USGS:15302200:00011:00014",
  "USGS:15302200:00011:00016",
  "USGS:15302200:00011:00003",
  "USGS:15302200:00011:00001",
  "USGS:15302200:00011:00013",
  "USGS:15302250:00011:00013",
  "USGS:15302250:00011:00015",
  "USGS:15302250:00011:00003",
  "USGS:15302250:00011:00001",
  "USGS:15302250:00011:00002",
  "USGS:15303900:00011:00002",
  "USGS:15303900:00011:00001",
  "USGS:15304000:00011:00016",
  "USGS:15304000:00011:00002",
  "USGS:15304000:00011:00003",
  "USGS:15304010:00011:00001",
  "USGS:15304010:00011:00002",
  "USGS:15320100:00011:00002",
  "USGS:15320100:00011:00001",
  "USGS:15348000:00011:00017",
  "USGS:15348000:00011:00001",
  "USGS:15348000:00011:00002",
  "USGS:15356000:00011:00003",
  "USGS:15356000:00011:00006",
  "USGS:15453500:00011:00017",
  "USGS:15453500:00011:00001",
  "USGS:15453500:00011:00003",
  "USGS:15457790:00011:00004",
  "USGS:15457790:00011:00001",
  "USGS:15457790:00011:00002",
  "USGS:15457800:00011:00001",
  "USGS:15457800:00011:00004",
  "USGS:15457800:00011:00002",
  "USGS:15457800:00011:00003",
  "USGS:15477740:00011:00015",
  "USGS:15477740:00011:00005",
  "USGS:15477740:00011:00002",
  "USGS:15477740:00011:00001",
  "USGS:15478038:00011:00002",
  "USGS:15478038:00011:00004",
  "USGS:15478038:00011:00014",
  "USGS:15478038:00011:00016",
  "USGS:15478038:00011:00020",
  "USGS:15478038:00011:00025",
  "USGS:15478038:00011:00019",
  "USGS:15478038:00011:00001",
  "USGS:15478038:00011:00023",
  "USGS:15478040:00011:00015",
  "USGS:15478040:00011:00016",
  "USGS:15478040:00011:00001",
  "USGS:15478040:00011:00002",
  "USGS:15484000:00011:00019",
  "USGS:15484000:00011:00015",
  "USGS:15484000:00011:00001",
  "USGS:15484000:00011:00002",
  "USGS:15485500:00011:00001",
  "USGS:15485500:00011:00002",
  "USGS:15493000:00011:00021",
  "USGS:15493000:00011:00022",
  "USGS:15493000:00011:00009",
  "USGS:15493000:00011:00001",
  "USGS:15493000:00011:00007",
  "USGS:15493000:00011:00023",
  "USGS:15502000:00011:00012",
  "USGS:15502000:00011:00014",
  "USGS:15502000:00011:00001",
  "USGS:15511000:00011:00020",
  "USGS:15511000:00011:00019",
  "USGS:15511000:00011:00002",
  "USGS:15511000:00011:00006",
  "USGS:15514000:00011:00002",
  "USGS:15514000:00011:00003",
  "USGS:15515060:00011:00003",
  "USGS:15515060:00011:00005",
  "USGS:15515060:00011:00001",
  "USGS:15515060:00011:00002",
  "USGS:15515500:00011:00001",
  "USGS:15515500:00011:00002",
  "USGS:15515500:00011:00003",
  "USGS:15519100:00011:00003",
  "USGS:15519100:00011:00014",
  "USGS:15519100:00011:00001",
  "USGS:15519100:00011:00002",
  "USGS:15519150:00011:00001",
  "USGS:15519150:00011:00002",
  "USGS:15564879:00011:00004",
  "USGS:15564879:00011:00002",
  "USGS:15564879:00011:00003",
  "USGS:15565447:00011:00001",
  "USGS:15565447:00011:00015",
  "USGS:15565447:00011:00002",
  "USGS:15565447:00011:00003",
  "USGS:15580095:00011:00003",
  "USGS:15580095:00011:00004",
  "USGS:15580095:00011:00002",
  "USGS:15580095:00011:00001",
  "USGS:15742980:00011:00002",
  "USGS:15743850:00011:00005",
  "USGS:15743850:00011:00017",
  "USGS:15743850:00011:00002",
  "USGS:15743850:00011:00001",
  "USGS:15744500:00011:00005",
  "USGS:15744500:00011:00006",
  "USGS:15747000:00011:00014",
  "USGS:15747000:00011:00015",
  "USGS:15747000:00011:00004",
  "USGS:15747000:00011:00002",
  "USGS:15803000:00011:00003",
  "USGS:15803000:00011:00004",
  "USGS:15803000:00011:00016",
  "USGS:15803000:00011:00001",
  "USGS:15803000:00011:00002",
  "USGS:15803000:00011:00014",
  "USGS:15820000:00011:00002",
  "USGS:15820000:00011:00014",
  "USGS:15875000:00011:00014",
  "USGS:15875000:00011:00004",
  "USGS:15875000:00011:00001",
  "USGS:15875000:00011:00015",
  "USGS:15875000:00011:00017",
  "USGS:15896000:00011:00001",
  "USGS:15896000:00011:00002",
  "USGS:15896000:00011:00003",
  "USGS:15905100:00011:00004",
  "USGS:15905100:00011:00003",
  "USGS:15905100:00011:00001",
  "USGS:15905100:00011:00002",
  "USGS:15908000:00011:00018",
  "USGS:15908000:00011:00015",
  "USGS:15908000:00011:00014",
  "USGS:15908000:00011:00001",
  "USGS:15908000:00011:00003",
  "USGS:15980000:00011:00004",
  "USGS:15980000:00011:00005",
  "USGS:15980000:00011:00001",
  "USGS:15980000:00011:00002",
  "USGS:16010000:00011:00001",
  "USGS:16010000:00011:00002",
  "USGS:611725149335401:00011:00001",
  "USGS:644528147131202:00011:00001",
  "USGS:644528147131202:00011:00003",
  "USGS:02197020:00011:00003",
  "USGS:02197020:00011:00002",
  "USGS:02197020:00011:00001",
  "USGS:021973269:00011:00003",
  "USGS:021973269:00011:00002",
  "USGS:021973269:00011:00001",
  "USGS:02197500:00011:00001",
  "USGS:02197500:00011:00003",
  "USGS:02197500:00011:00002",
  "USGS:02197598:00011:00002",
  "USGS:02197598:00011:00001",
  "USGS:02197830:00011:00003",
  "USGS:02197830:00011:00001",
  "USGS:02197830:00011:00002",
  "USGS:02198000:00011:00007",
  "USGS:02198000:00011:00002",
  "USGS:02198000:00011:00003",
  "USGS:02198100:00011:00003",
  "USGS:02198100:00011:00001",
  "USGS:02198100:00011:00002",
  "USGS:02198375:00011:00003",
  "USGS:02198375:00011:00001",
  "USGS:02198500:00011:00001",
  "USGS:02198500:00011:00002",
  "USGS:02198690:00011:00002",
  "USGS:02198690:00011:00001",
  "USGS:02198759:00011:00005",
  "USGS:02198759:00011:00007",
  "USGS:02198759:00011:00002",
  "USGS:02198759:00011:00001",
  "USGS:02198810:00011:00019",
  "USGS:02198810:00011:00004",
  "USGS:02198810:00011:00005",
  "USGS:02198810:00011:00018",
  "USGS:02198810:00011:00003",
  "USGS:02198810:00011:00020",
  "USGS:02198810:00011:00034",
  "USGS:02198810:00011:00033",
  "USGS:02198810:00011:00035",
  "USGS:02198820:00011:00004",
  "USGS:02198820:00011:00011",
  "USGS:02198820:00011:00013",
  "USGS:02198820:00011:00010",
  "USGS:02198820:00011:00009",
  "USGS:02198820:00011:00002",
  "USGS:02198820:00011:00012",
  "USGS:02198820:00011:00001",
  "USGS:02198820:00011:00005",
  "USGS:02198820:00011:00006",
  "USGS:02198820:00011:00008",
  "USGS:02198820:00011:00007",
  "USGS:02198840:00011:00013",
  "USGS:02198840:00011:00004",
  "USGS:02198840:00011:00023",
  "USGS:02198840:00011:00003",
  "USGS:02198840:00011:00002",
  "USGS:02198840:00011:00020",
  "USGS:02198840:00011:00021",
  "USGS:02198840:00011:00018",
  "USGS:02198840:00011:00022",
  "USGS:02198920:00011:00006",
  "USGS:02198920:00011:00012",
  "USGS:02198920:00011:00023",
  "USGS:02198920:00011:00027",
  "USGS:02198920:00011:00001",
  "USGS:02198920:00011:00004",
  "USGS:02198920:00011:00022",
  "USGS:02198920:00011:00041",
  "USGS:02198920:00011:00021",
  "USGS:02198920:00011:00042",
  "USGS:02198950:00011:00029",
  "USGS:02198950:00011:00002",
  "USGS:02198950:00011:00015",
  "USGS:02198950:00011:00001",
  "USGS:02198950:00011:00030",
  "USGS:02198950:00011:00031",
  "USGS:02198950:00011:00032",
  "USGS:02198950:00011:00033",
  "USGS:02198955:00011:00009",
  "USGS:02198955:00011:00004",
  "USGS:02198955:00011:00005",
  "USGS:02198955:00011:00001",
  "USGS:02198955:00011:00010",
  "USGS:02198955:00011:00013",
  "USGS:02198955:00011:00011",
  "USGS:02198955:00011:00012",
  "USGS:021989715:00011:00001",
  "USGS:021989715:00011:00006",
  "USGS:021989715:00011:00021",
  "USGS:021989715:00011:00002",
  "USGS:021989715:00011:00007",
  "USGS:021989715:00011:00003",
  "USGS:021989715:00011:00018",
  "USGS:021989715:00011:00004",
  "USGS:021989715:00011:00005",
  "USGS:021989715:00011:00019",
  "USGS:021989715:00011:00017",
  "USGS:021989715:00011:00020",
  "USGS:021989773:00011:00007",
  "USGS:021989773:00011:00014",
  "USGS:021989773:00011:00015",
  "USGS:021989773:00011:00012",
  "USGS:021989773:00011:00011",
  "USGS:021989773:00011:00002",
  "USGS:021989773:00011:00003",
  "USGS:021989773:00011:00025",
  "USGS:021989773:00011:00001",
  "USGS:021989773:00011:00008",
  "USGS:021989773:00011:00009",
  "USGS:021989773:00011:00010",
  "USGS:021989773:00011:00026",
  "USGS:021989773:00011:00042",
  "USGS:021989792:00011:00029",
  "USGS:021989792:00011:00002",
  "USGS:021989792:00011:00015",
  "USGS:021989792:00011:00001",
  "USGS:021989792:00011:00030",
  "USGS:021989792:00011:00031",
  "USGS:021989792:00011:00032",
  "USGS:021989792:00011:00033",
  "USGS:021989793:00011:00001",
  "USGS:021989793:00011:00002",
  "USGS:021989793:00011:00005",
  "USGS:021989793:00011:00003",
  "USGS:021989793:00011:00004",
  "USGS:0219897945:00011:00001",
  "USGS:0219897945:00011:00002",
  "USGS:0219897945:00011:00005",
  "USGS:0219897945:00011:00003",
  "USGS:0219897945:00011:00004",
  "USGS:02198980:00011:00036",
  "USGS:02198980:00011:00004",
  "USGS:02198980:00011:00005",
  "USGS:02198980:00011:00003",
  "USGS:02198980:00011:00008",
  "USGS:02198980:00011:00022",
  "USGS:02198980:00011:00001",
  "USGS:02198980:00011:00037",
  "USGS:02199000:00011:00006",
  "USGS:02199000:00011:00007",
  "USGS:02199000:00011:00003",
  "USGS:02199000:00011:00002",
  "USGS:02199000:00011:00005",
  "USGS:02199000:00011:00001",
  "USGS:02200120:00011:00005",
  "USGS:02200120:00011:00004",
  "USGS:02200120:00011:00003",
  "USGS:02201000:00011:00016",
  "USGS:02201000:00011:00001",
  "USGS:02201000:00011:00002",
  "USGS:02201230:00011:00003",
  "USGS:02201230:00011:00002",
  "USGS:02201230:00011:00001",
  "USGS:02202040:00011:00002",
  "USGS:02202040:00011:00007",
  "USGS:02202040:00011:00001",
  "USGS:02202190:00011:00005",
  "USGS:02202190:00011:00004",
  "USGS:02202190:00011:00003",
  "USGS:02202500:00011:00002",
  "USGS:02202500:00011:00006",
  "USGS:02202600:00011:00003",
  "USGS:02202600:00011:00001",
  "USGS:02202600:00011:00002",
  "USGS:02202680:00011:00003",
  "USGS:02202680:00011:00002",
  "USGS:02202680:00011:00001",
  "USGS:02203000:00011:00001",
  "USGS:02203000:00011:00002",
  "USGS:02203518:00011:00003",
  "USGS:02203518:00011:00001",
  "USGS:02203518:00011:00002",
  "USGS:02203536:00011:00023",
  "USGS:02203536:00011:00003",
  "USGS:02203536:00011:00004",
  "USGS:02203536:00011:00002",
  "USGS:02203536:00011:00001",
  "USGS:02203559:00011:00003",
  "USGS:02203559:00011:00001",
  "USGS:02203559:00011:00002",
  "USGS:022035975:00011:00003",
  "USGS:022035975:00011:00012",
  "USGS:022035975:00011:00036",
  "USGS:022035975:00011:00009",
  "USGS:022035975:00011:00010",
  "USGS:022035975:00011:00002",
  "USGS:022035975:00011:00001",
  "USGS:022035975:00011:00004",
  "USGS:022035975:00011:00006",
  "USGS:022035975:00011:00007",
  "USGS:022035975:00011:00037",
  "USGS:022035975:00011:00008",
  "USGS:02203603:00011:00013",
  "USGS:02203603:00011:00003",
  "USGS:02203603:00011:00002",
  "USGS:02203603:00011:00001",
  "USGS:02203603:00011:00014",
  "USGS:02203603:00011:00015",
  "USGS:02203603:00011:00016",
  "USGS:02203603:00011:00017",
  "USGS:02203655:00011:00004",
  "USGS:02203655:00011:00003",
  "USGS:02203655:00011:00002",
  "USGS:02203655:00011:00001",
  "USGS:02203655:00011:00005",
  "USGS:02203655:00011:00006",
  "USGS:02203655:00011:00007",
  "USGS:02203655:00011:00008",
  "USGS:02203700:00011:00011",
  "USGS:02203700:00011:00005",
  "USGS:02203700:00011:00004",
  "USGS:02207135:00011:00010",
  "USGS:02203700:00011:00003",
  "USGS:02203700:00011:00006",
  "USGS:02203700:00011:00007",
  "USGS:02203700:00011:00008",
  "USGS:02203700:00011:00009",
  "USGS:02203831:00011:00016",
  "USGS:02203831:00011:00006",
  "USGS:02203831:00011:00003",
  "USGS:02203831:00011:00017",
  "USGS:02203831:00011:00018",
  "USGS:02203831:00011:00019",
  "USGS:02203831:00011:00020",
  "USGS:02203863:00011:00014",
  "USGS:02203863:00011:00003",
  "USGS:02203863:00011:00002",
  "USGS:02203863:00011:00001",
  "USGS:02203863:00011:00015",
  "USGS:02203863:00011:00018",
  "USGS:02203863:00011:00016",
  "USGS:02203863:00011:00017",
  "USGS:02203873:00011:00007",
  "USGS:02203873:00011:00005",
  "USGS:02203873:00011:00004",
  "USGS:02203873:00011:00008",
  "USGS:02203873:00011:00010",
  "USGS:02203873:00011:00009",
  "USGS:02203873:00011:00011",
  "USGS:02203900:00011:00008",
  "USGS:02203900:00011:00007",
  "USGS:02203900:00011:00004",
  "USGS:02203900:00011:00003",
  "USGS:02203900:00011:00009",
  "USGS:02203900:00011:00012",
  "USGS:02203900:00011:00010",
  "USGS:02203900:00011:00011",
  "USGS:02203950:00011:00014",
  "USGS:02203950:00011:00003",
  "USGS:02203950:00011:00002",
  "USGS:02203950:00011:00001",
  "USGS:02203950:00011:00015",
  "USGS:02203950:00011:00016",
  "USGS:02203950:00011:00017",
  "USGS:02203950:00011:00018",
  "USGS:02203960:00011:00014",
  "USGS:02203960:00011:00004",
  "USGS:02203960:00011:00002",
  "USGS:02203960:00011:00001",
  "USGS:02203960:00011:00015",
  "USGS:02203960:00011:00016",
  "USGS:02203960:00011:00017",
  "USGS:02203960:00011:00018",
  "USGS:02204037:00011:00005",
  "USGS:02204037:00011:00003",
  "USGS:02204037:00011:00002",
  "USGS:02204037:00011:00006",
  "USGS:02204037:00011:00010",
  "USGS:02204037:00011:00007",
  "USGS:02204037:00011:00008",
  "USGS:02204070:00011:00008",
  "USGS:02204070:00011:00002",
  "USGS:02204070:00011:00004",
  "USGS:02204130:00011:00003",
  "USGS:02204130:00011:00002",
  "USGS:02204130:00011:00001",
  "USGS:02204285:00011:00003",
  "USGS:02204285:00011:00001",
  "USGS:02204285:00011:00002",
  "USGS:09379200:00011:00015",
  "USGS:09379200:00011:00004",
  "USGS:09379200:00011:00003",
  "USGS:09380000:00011:00003",
  "USGS:09380000:00011:00014",
  "USGS:09380000:00011:00001",
  "USGS:09380000:00011:00002",
  "USGS:09380000:00011:00004",
  "USGS:09382000:00011:00001",
  "USGS:09382000:00011:00002",
  "USGS:09383300:00011:00001",
  "USGS:09383300:00011:00002",
  "USGS:09383400:00011:00015",
  "USGS:09383400:00011:00001",
  "USGS:09383400:00011:00002",
  "USGS:09383409:00011:00004",
  "USGS:09383409:00011:00001",
  "USGS:09383409:00011:00003",
  "USGS:09383417:00011:00004",
  "USGS:09383417:00011:00001",
  "USGS:09383417:00011:00003",
  "USGS:09383500:00011:00015",
  "USGS:02207135:00011:00011",
  "USGS:02207160:00011:00005",
  "USGS:02207160:00011:00003",
  "USGS:02207160:00011:00002",
  "USGS:02207160:00011:00006",
  "USGS:02207160:00011:00009",
  "USGS:02207160:00011:00007",
  "USGS:02207160:00011:00008",
  "USGS:02207185:00011:00004",
  "USGS:02207185:00011:00003",
  "USGS:02207185:00011:00002",
  "USGS:02207185:00011:00001",
  "USGS:02207185:00011:00005",
  "USGS:02207200:00011:00004",
  "USGS:02207200:00011:00003",
  "USGS:02207220:00011:00003",
  "USGS:02207220:00011:00002",
  "USGS:02207220:00011:00001",
  "USGS:02207300:00011:00008",
  "USGS:02207300:00011:00007",
  "USGS:02207335:00011:00006",
  "USGS:02207335:00011:00002",
  "USGS:02207335:00011:00001",
  "USGS:02207385:00011:00004",
  "USGS:02207385:00011:00003",
  "USGS:02207385:00011:00002",
  "USGS:02207385:00011:00001",
  "USGS:02207385:00011:00006",
  "USGS:02207400:00011:00004",
  "USGS:02207400:00011:00003",
  "USGS:02207400:00011:00002",
  "USGS:02207400:00011:00001",
  "USGS:02207400:00011:00006",
  "USGS:02207414:00011:00006",
  "USGS:02207414:00011:00008",
  "USGS:02207414:00011:00005",
  "USGS:02207414:00011:00004",
  "USGS:02207414:00011:00002",
  "USGS:02207414:00011:00007",
  "USGS:02207414:00011:00001",
  "USGS:02207418:00011:00002",
  "USGS:02207418:00011:00017",
  "USGS:02207418:00011:00001",
  "USGS:02207435:00011:00002",
  "USGS:02207435:00011:00004",
  "USGS:02207435:00011:00001",
  "USGS:02207448:00011:00003",
  "USGS:02207448:00011:00015",
  "USGS:02207448:00011:00002",
  "USGS:02207448:00011:00001",
  "USGS:02208000:00011:00003",
  "USGS:02208000:00011:00002",
  "USGS:02208000:00011:00001",
  "USGS:02208050:00011:00002",
  "USGS:02208050:00011:00003",
  "USGS:02208050:00011:00001",
  "USGS:02208150:00011:00004",
  "USGS:02352500:00011:00001",
  "USGS:02208150:00011:00003",
  "USGS:02208150:00011:00002",
  "USGS:02208150:00011:00001",
  "USGS:02208150:00011:00007",
  "USGS:02208450:00011:00015",
  "USGS:02208450:00011:00004",
  "USGS:02208450:00011:00002",
  "USGS:02208450:00011:00003",
  "USGS:02208450:00011:00016",
  "USGS:02208450:00011:00019",
  "USGS:02208450:00011:00017",
  "USGS:02208450:00011:00018",
  "USGS:02208485:00011:00004",
  "USGS:02208485:00011:00001",
  "USGS:02208487:00011:00001",
  "USGS:02208493:00011:00014",
  "USGS:02208493:00011:00003",
  "USGS:02208493:00011:00002",
  "USGS:02208493:00011:00001",
  "USGS:02208493:00011:00015",
  "USGS:02208493:00011:00018",
  "USGS:02208493:00011:00016",
  "USGS:02208493:00011:00017",
  "USGS:02209000:00011:00003",
  "USGS:02209000:00011:00001",
  "USGS:02209000:00011:00002",
  "USGS:02209360:00011:00003",
  "USGS:02209360:00011:00002",
  "USGS:02209360:00011:00001",
  "USGS:02210500:00011:00001",
  "USGS:02210500:00011:00002",
  "USGS:02211375:00011:00003",
  "USGS:02211375:00011:00002",
  "USGS:02211375:00011:00001",
  "USGS:02211800:00011:00004",
  "USGS:02211800:00011:00005",
  "USGS:02211800:00011:00003",
  "USGS:02212600:00011:00001",
  "USGS:02212600:00011:00002",
  "USGS:02212600:00011:00003",
  "USGS:02212735:00011:00003",
  "USGS:02212735:00011:00001",
  "USGS:02212735:00011:00002",
  "USGS:02213000:00011:00009",
  "USGS:02213000:00011:00002",
  "USGS:02213000:00011:00006",
  "USGS:02213500:00011:00005",
  "USGS:02213500:00011:00001",
  "USGS:02213500:00011:00002",
  "USGS:02214075:00011:00003",
  "USGS:02214075:00011:00002",
  "USGS:02214075:00011:00001",
  "USGS:02214590:00011:00003",
  "USGS:02214590:00011:00001",
  "USGS:02214590:00011:00002",
  "USGS:02215000:00011:00014",
  "USGS:02215000:00011:00003",
  "USGS:02215000:00011:00001",
  "USGS:02215000:00011:00002",
  "USGS:02215100:00011:00001",
  "USGS:02215100:00011:00002",
  "USGS:02215260:00011:00016",
  "USGS:02215260:00011:00005",
  "USGS:02215260:00011:00002",
  "USGS:02215260:00011:00001",
  "USGS:02215500:00011:00001",
  "USGS:02215500:00011:00006",
  "USGS:02215500:00011:00002",
  "USGS:02215500:00011:00003",
  "USGS:02215900:00011:00003",
  "USGS:02215900:00011:00002",
  "USGS:02215900:00011:00001",
  "USGS:02216180:00011:00003",
  "USGS:02216180:00011:00001",
  "USGS:02216180:00011:00002",
  "USGS:02217274:00011:00004",
  "USGS:02217274:00011:00003",
  "USGS:02217274:00011:00002",
  "USGS:02217274:00011:00001",
  "USGS:02217274:00011:00005",
  "USGS:02217297:00011:00003",
  "USGS:02217297:00011:00002",
  "USGS:02217297:00011:00001",
  "USGS:02217475:00011:00005",
  "USGS:02217475:00011:00001",
  "USGS:02217475:00011:00002",
  "USGS:02217500:00011:00001",
  "USGS:02217500:00011:00002",
  "USGS:02217615:00011:00003",
  "USGS:02217615:00011:00002",
  "USGS:02217615:00011:00001",
  "USGS:02217643:00011:00005",
  "USGS:02217643:00011:00004",
  "USGS:02217643:00011:00001",
  "USGS:02217643:00011:00006",
  "USGS:02217643:00011:00007",
  "USGS:02217643:00011:00008",
  "USGS:02217643:00011:00009",
  "USGS:02217770:00011:00003",
  "USGS:02217770:00011:00002",
  "USGS:02217770:00011:00001",
  "USGS:02381400:00011:00006",
  "USGS:02381400:00011:00007",
  "USGS:02381400:00011:00004",
  "USGS:02381400:00011:00003",
  "USGS:02381400:00011:00002",
  "USGS:02381400:00011:00001",
  "USGS:02381400:00011:00017",
  "USGS:09482000:00011:00001",
  "USGS:09482000:00011:00002",
  "USGS:09482500:00011:00003",
  "USGS:09482500:00011:00004",
  "USGS:09484000:00011:00003",
  "USGS:09484000:00011:00001",
  "USGS:09484000:00011:00002",
  "USGS:09484500:00011:00001",
  "USGS:09484500:00011:00002",
  "USGS:09484550:00011:00003",
  "USGS:09484550:00011:00001",
  "USGS:02338500:00011:00024",
  "USGS:02338500:00011:00007",
  "USGS:02338500:00011:00009",
  "USGS:02338500:00011:00001",
  "USGS:02338500:00011:00006",
  "USGS:02338523:00011:00027",
  "USGS:02338523:00011:00003",
  "USGS:02338523:00011:00002",
  "USGS:02338523:00011:00001",
  "USGS:02338660:00011:00006",
  "USGS:02338660:00011:00002",
  "USGS:02338660:00011:00003",
  "USGS:02338840:00011:00013",
  "USGS:02338840:00011:00002",
  "USGS:02338840:00011:00003",
  "USGS:02339400:00011:00006",
  "USGS:02339400:00011:00007",
  "USGS:02339400:00011:00004",
  "USGS:02339400:00011:00003",
  "USGS:02339400:00011:00002",
  "USGS:02339400:00011:00001",
  "USGS:02339400:00011:00018",
  "USGS:02339402:00011:00001",
  "USGS:02339500:00011:00005",
  "USGS:02339500:00011:00001",
  "USGS:02339500:00011:00002",
  "USGS:02341460:00011:00005",
  "USGS:02341460:00011:00006",
  "USGS:02341460:00011:00009",
  "USGS:02341460:00011:00008",
  "USGS:02341460:00011:00004",
  "USGS:02341460:00011:00007",
  "USGS:02341460:00011:00002",
  "USGS:02341460:00011:00001",
  "USGS:02341505:00011:00003",
  "USGS:02341505:00011:00006",
  "USGS:02341505:00011:00001",
  "USGS:02341800:00011:00013",
  "USGS:02341800:00011:00001",
  "USGS:02341800:00011:00002",
  "USGS:02342850:00011:00005",
  "USGS:02342850:00011:00001",
  "USGS:02342850:00011:00004",
  "USGS:02342881:00011:00004",
  "USGS:02342881:00011:00005",
  "USGS:02342881:00011:00003",
  "USGS:02343225:00011:00005",
  "USGS:02343225:00011:00004",
  "USGS:02343225:00011:00003",
  "USGS:02343240:00011:00006",
  "USGS:02343240:00011:00007",
  "USGS:02343240:00011:00004",
  "USGS:02343240:00011:00003",
  "USGS:02343240:00011:00002",
  "USGS:02343240:00011:00001",
  "USGS:02343240:00011:00017",
  "USGS:02343241:00011:00001",
  "USGS:02343801:00011:00032",
  "USGS:02343801:00011:00033",
  "USGS:02343801:00011:00020",
  "USGS:02343801:00011:00013",
  "USGS:02343801:00011:00014",
  "USGS:02343801:00011:00015",
  "USGS:02343801:00011:00016",
  "USGS:02343801:00011:00017",
  "USGS:02343801:00011:00018",
  "USGS:02343801:00011:00035",
  "USGS:02343805:00011:00013",
  "USGS:02343805:00011:00001",
  "USGS:02343805:00011:00002",
  "USGS:02343940:00011:00002",
  "USGS:02343940:00011:00004",
  "USGS:02343940:00011:00001",
  "USGS:02344280:00011:00014",
  "USGS:02344280:00011:00004",
  "USGS:02344280:00011:00001",
  "USGS:02344327:00011:00004",
  "USGS:02344327:00011:00001",
  "USGS:02344350:00011:00003",
  "USGS:02344350:00011:00001",
  "USGS:02344350:00011:00002",
  "USGS:02344396:00011:00003",
  "USGS:02344396:00011:00002",
  "USGS:02344396:00011:00001",
  "USGS:02344423:00011:00006",
  "USGS:02344423:00011:00008",
  "USGS:02344423:00011:00005",
  "USGS:02344423:00011:00004",
  "USGS:02344423:00011:00003",
  "USGS:02344423:00011:00007",
  "USGS:02344423:00011:00001",
  "USGS:02344424:00011:00001",
  "USGS:02344478:00011:00004",
  "USGS:02344478:00011:00001",
  "USGS:02344478:00011:00002",
  "USGS:02344500:00011:00001",
  "USGS:02344500:00011:00002",
  "USGS:02344605:00011:00002",
  "USGS:02344605:00011:00001",
  "USGS:02344620:00011:00002",
  "USGS:02344620:00011:00003",
  "USGS:02344620:00011:00001",
  "USGS:02344630:00011:00004",
  "USGS:02344630:00011:00003",
  "USGS:02344630:00011:00002",
  "USGS:02344630:00011:00001",
  "USGS:02344630:00011:00005",
  "USGS:02344630:00011:00006",
  "USGS:02344630:00011:00007",
  "USGS:02344630:00011:00008",
  "USGS:02344650:00011:00007",
  "USGS:02344650:00011:00009",
  "USGS:02344650:00011:00006",
  "USGS:02344650:00011:00005",
  "USGS:02344650:00011:00004",
  "USGS:02344650:00011:00008",
  "USGS:02344650:00011:00001",
  "USGS:02344655:00011:00003",
  "USGS:02344655:00011:00002",
  "USGS:02344655:00011:00001",
  "USGS:02344655:00011:00004",
  "USGS:02344655:00011:00005",
  "USGS:02344671:00011:00006",
  "USGS:02344671:00011:00008",
  "USGS:02344671:00011:00005",
  "USGS:02344671:00011:00004",
  "USGS:02344671:00011:00003",
  "USGS:02344671:00011:00007",
  "USGS:02344671:00011:00001",
  "USGS:02344673:00011:00003",
  "USGS:02344673:00011:00001",
  "USGS:02344673:00011:00004",
  "USGS:02344673:00011:00007",
  "USGS:02344673:00011:00005",
  "USGS:02344673:00011:00006",
  "USGS:02344700:00011:00001",
  "USGS:02344700:00011:00002",
  "USGS:02344724:00011:00004",
  "USGS:02344724:00011:00001",
  "USGS:02344736:00011:00004",
  "USGS:02344736:00011:00001",
  "USGS:02344748:00011:00004",
  "USGS:02344748:00011:00001",
  "USGS:02344872:00011:00003",
  "USGS:02344872:00011:00002",
  "USGS:02344872:00011:00001",
  "USGS:02346310:00011:00003",
  "USGS:02346310:00011:00002",
  "USGS:02346310:00011:00001",
  "USGS:02347500:00011:00007",
  "USGS:02347500:00011:00002",
  "USGS:02347500:00011:00006",
  "USGS:02349605:00011:00003",
  "USGS:02349605:00011:00001",
  "USGS:02349605:00011:00002",
  "USGS:02349900:00011:00003",
  "USGS:02349900:00011:00001",
  "USGS:02349900:00011:00002",
  "USGS:02350512:00011:00006",
  "USGS:02350512:00011:00001",
  "USGS:02350512:00011:00002",
  "USGS:02350600:00011:00005",
  "USGS:02350600:00011:00001",
  "USGS:02350600:00011:00002",
  "USGS:02350900:00011:00009",
  "USGS:02350900:00011:00005",
  "USGS:02350900:00011:00001",
  "USGS:02350900:00011:00002",
  "USGS:02351500:00011:00003",
  "USGS:02351500:00011:00002",
  "USGS:02351500:00011:00001",
  "USGS:02351890:00011:00005",
  "USGS:02351890:00011:00001",
  "USGS:02351890:00011:00002",
  "USGS:02352500:00011:00008",
  "USGS:02352500:00011:00002",
  "USGS:02352500:00011:00003",
  "USGS:02352500:00011:00009",
  "USGS:02353000:00011:00023",
  "USGS:02353000:00011:00006",
  "USGS:02353000:00011:00001",
  "USGS:02353000:00011:00002",
  "USGS:07381331:00011:00003",
  "USGS:07381331:00011:00002",
  "USGS:07381331:00011:00004",
  "USGS:07381331:00011:00016",
  "USGS:07381331:00011:00014",
  "USGS:07381331:00011:00017",
  "USGS:07381331:00011:00018",
  "USGS:09507580:00011:00003",
  "USGS:09507580:00011:00001",
  "USGS:09507580:00011:00002",
  "USGS:09507980:00011:00003",
  "USGS:09507980:00011:00001",
  "USGS:09507980:00011:00002",
  "USGS:09508000:00011:00003",
  "USGS:09508000:00011:00002",
  "USGS:09508300:00011:00004",
  "USGS:09508300:00011:00003",
  "USGS:09508500:00011:00003",
  "USGS:09508500:00011:00005",
  "USGS:09508500:00011:00006",
  "USGS:09509501:00011:00001",
  "USGS:09509501:00011:00003",
  "USGS:02218300:00011:00005",
  "USGS:02218300:00011:00001",
  "USGS:02218300:00011:00002",
  "USGS:02218565:00011:00004",
  "USGS:02218565:00011:00003",
  "USGS:02218565:00011:00002",
  "USGS:02218565:00011:00001",
  "USGS:02218565:00011:00005",
  "USGS:02219000:00011:00018",
  "USGS:02219000:00011:00001",
  "USGS:02219000:00011:00002",
  "USGS:02220788:00011:00002",
  "USGS:02220788:00011:00001",
  "USGS:02220900:00011:00008",
  "USGS:02220900:00011:00001",
  "USGS:02220900:00011:00002",
  "USGS:02221525:00011:00001",
  "USGS:02221525:00011:00002",
  "USGS:02223000:00011:00008",
  "USGS:02223000:00011:00002",
  "USGS:02223000:00011:00003",
  "USGS:02223056:00011:00020",
  "USGS:02223056:00011:00008",
  "USGS:02223056:00011:00002",
  "USGS:02223056:00011:00001",
  "USGS:02223110:00011:00013",
  "USGS:02223110:00011:00002",
  "USGS:02223110:00011:00001",
  "USGS:02223190:00011:00002",
  "USGS:02223190:00011:00012",
  "USGS:02223190:00011:00001",
  "USGS:02223248:00011:00002",
  "USGS:02223248:00011:00001",
  "USGS:02223360:00011:00003",
  "USGS:02223360:00011:00001",
  "USGS:02223360:00011:00002",
  "USGS:02223500:00011:00010",
  "USGS:02223500:00011:00002",
  "USGS:02223500:00011:00006",
  "USGS:02224500:00011:00005",
  "USGS:02224500:00011:00001",
  "USGS:02224500:00011:00002",
  "USGS:02224940:00011:00014",
  "USGS:02224940:00011:00003",
  "USGS:02224940:00011:00002",
  "USGS:02224940:00011:00001",
  "USGS:02225000:00011:00001",
  "USGS:02225000:00011:00013",
  "USGS:02225000:00011:00002",
  "USGS:02225000:00011:00003",
  "USGS:02225270:00011:00005",
  "USGS:02225270:00011:00004",
  "USGS:02225270:00011:00003",
  "USGS:02225500:00011:00007",
  "USGS:02225500:00011:00002",
  "USGS:02225500:00011:00003",
  "USGS:02226000:00011:00001",
  "USGS:02226000:00011:00010",
  "USGS:02226000:00011:00002",
  "USGS:02226000:00011:00003",
  "USGS:02226160:00011:00025",
  "USGS:02226160:00011:00010",
  "USGS:02226160:00011:00008",
  "USGS:02226160:00011:00007",
  "USGS:022261794:00011:00006",
  "USGS:022261794:00011:00007",
  "USGS:022261794:00011:00002",
  "USGS:022261794:00011:00001",
  "USGS:02226180:00011:00003",
  "USGS:02226180:00011:00004",
  "USGS:02226180:00011:00002",
  "USGS:02226180:00011:00001",
  "USGS:02226362:00011:00003",
  "USGS:02226362:00011:00001",
  "USGS:02226362:00011:00002",
  "USGS:02226500:00011:00001",
  "USGS:02226500:00011:00006",
  "USGS:02226500:00011:00002",
  "USGS:02226500:00011:00003",
  "USGS:02227270:00011:00002",
  "USGS:02227270:00011:00012",
  "USGS:02227270:00011:00001",
  "USGS:02227500:00011:00003",
  "USGS:02227500:00011:00001",
  "USGS:02227500:00011:00002",
  "USGS:02228000:00011:00001",
  "USGS:02228000:00011:00008",
  "USGS:02228000:00011:00002",
  "USGS:02228000:00011:00004",
  "USGS:02228070:00011:00018",
  "USGS:02228070:00011:00003",
  "USGS:02228070:00011:00013",
  "USGS:02228070:00011:00001",
  "USGS:02228070:00011:00002",
  "USGS:02228295:00011:00010",
  "USGS:02228295:00011:00011",
  "USGS:02228295:00011:00009",
  "USGS:02228295:00011:00008",
  "USGS:02228295:00011:00002",
  "USGS:02228295:00011:00001",
  "USGS:02231254:00011:00018",
  "USGS:02231254:00011:00007",
  "USGS:02231254:00011:00003",
  "USGS:02231254:00011:00002",
  "USGS:02231254:00011:00001",
  "USGS:02314495:00011:00002",
  "USGS:02314495:00011:00001",
  "USGS:02314500:00011:00010",
  "USGS:02314500:00011:00007",
  "USGS:02314500:00011:00001",
  "USGS:02314500:00011:00002",
  "USGS:02315920:00011:00003",
  "USGS:02315920:00011:00001",
  "USGS:02315920:00011:00002",
  "USGS:02316000:00011:00004",
  "USGS:02316000:00011:00002",
  "USGS:02316000:00011:00003",
  "USGS:02317500:00011:00001",
  "USGS:02317500:00011:00027",
  "USGS:02317500:00011:00021",
  "USGS:02317500:00011:00022",
  "USGS:02317500:00011:00007",
  "USGS:02317500:00011:00026",
  "USGS:02317500:00011:00002",
  "USGS:02317500:00011:00006",
  "USGS:023177483:00011:00006",
  "USGS:023177483:00011:00002",
  "USGS:023177483:00011:00001",
  "USGS:02317755:00011:00004",
  "USGS:02317755:00011:00002",
  "USGS:02317797:00011:00014",
  "USGS:02317797:00011:00002",
  "USGS:02317797:00011:00003",
  "USGS:02317797:00011:00001",
  "USGS:02318000:00011:00003",
  "USGS:02318000:00011:00001",
  "USGS:02318000:00011:00002",
  "USGS:02318380:00011:00003",
  "USGS:02318380:00011:00002",
  "USGS:02318380:00011:00001",
  "USGS:02318500:00011:00006",
  "USGS:02318500:00011:00004",
  "USGS:02318500:00011:00001",
  "USGS:02318500:00011:00002",
  "USGS:02318700:00011:00015",
  "USGS:02318700:00011:00003",
  "USGS:02318700:00011:00001",
  "USGS:02318700:00011:00002",
  "USGS:02327355:00011:00003",
  "USGS:02327355:00011:00002",
  "USGS:02327355:00011:00001",
  "USGS:02327500:00011:00021",
  "USGS:02327500:00011:00017",
  "USGS:02327500:00011:00003",
  "USGS:02327500:00011:00001",
  "USGS:02327500:00011:00002",
  "USGS:02329342:00011:00003",
  "USGS:02329342:00011:00002",
  "USGS:02329342:00011:00001",
  "USGS:02330450:00011:00007",
  "USGS:02330450:00011:00008",
  "USGS:02330450:00011:00023",
  "USGS:02330450:00011:00021",
  "USGS:02330450:00011:00020",
  "USGS:02330450:00011:00005",
  "USGS:02330450:00011:00024",
  "USGS:02330450:00011:00001",
  "USGS:02330450:00011:00002",
  "USGS:02331000:00011:00005",
  "USGS:02331000:00011:00002",
  "USGS:02331000:00011:00004",
  "USGS:023312495:00011:00003",
  "USGS:023312495:00011:00002",
  "USGS:023312495:00011:00001",
  "USGS:02331600:00011:00003",
  "USGS:02331600:00011:00001",
  "USGS:02331600:00011:00002",
  "USGS:02381401:00011:00001",
  "USGS:02393377:00011:00002",
  "USGS:02393377:00011:00001",
  "USGS:02393419:00011:00003",
  "USGS:02393419:00011:00002",
  "USGS:02393419:00011:00001",
  "USGS:02393500:00011:00008",
  "USGS:02393500:00011:00009",
  "USGS:02393500:00011:00006",
  "USGS:02393500:00011:00005",
  "USGS:02393500:00011:00004",
  "USGS:02393500:00011:00002",
  "USGS:02393500:00011:00019",
  "USGS:02393501:00011:00001",
  "USGS:02394000:00011:00001",
  "USGS:02394000:00011:00002",
  "USGS:02394000:00011:00003",
  "USGS:02394670:00011:00016",
  "USGS:02394670:00011:00018",
  "USGS:02394670:00011:00001",
  "USGS:02394820:00011:00015",
  "USGS:02394820:00011:00003",
  "USGS:02394820:00011:00002",
  "USGS:02394820:00011:00001",
  "USGS:02395000:00011:00001",
  "USGS:02395000:00011:00002",
  "USGS:02395120:00011:00001",
  "USGS:02395120:00011:00002",
  "USGS:02395980:00011:00002",
  "USGS:02395980:00011:00001",
  "USGS:02395996:00011:00001",
  "USGS:02397000:00011:00001",
  "USGS:02397000:00011:00008",
  "USGS:02397000:00011:00002",
  "USGS:02397000:00011:00003",
  "USGS:02397410:00011:00005",
  "USGS:02397410:00011:00001",
  "USGS:02397410:00011:00002",
  "USGS:02397500:00011:00005",
  "USGS:02397500:00011:00001",
  "USGS:02397500:00011:00002",
  "USGS:02398000:00011:00001",
  "USGS:02398000:00011:00002",
  "USGS:02411930:00011:00002",
  "USGS:02411930:00011:00001",
  "USGS:02413000:00011:00005",
  "USGS:02413000:00011:00001",
  "USGS:02413000:00011:00004",
  "USGS:02413210:00011:00003",
  "USGS:02413210:00011:00002",
  "USGS:02413210:00011:00001",
  "USGS:03544970:00011:00014",
  "USGS:03544970:00011:00003",
  "USGS:03544970:00011:00002",
  "USGS:03544970:00011:00001",
  "USGS:03550500:00011:00014",
  "USGS:03550500:00011:00001",
  "USGS:03550500:00011:00002",
  "USGS:03567340:00011:00005",
  "USGS:03567340:00011:00004",
  "USGS:03567340:00011:00003",
  "USGS:03568933:00011:00005",
  "USGS:03568933:00011:00002",
  "USGS:03568933:00011:00003",
  "USGS:304406081330502:00011:00001",
  "USGS:304406081330503:00011:00001",
  "USGS:304406081330504:00011:00001",
  "USGS:304406081330505:00011:00001",
  "USGS:304949083165301:00011:00001",
  "USGS:305736084355801:00011:00001",
  "USGS:310507084262201:00011:00001",
  "USGS:310651084404501:00011:00001",
  "USGS:310810081292801:00011:00001",
  "USGS:310810081292802:00011:00002",
  "USGS:310810081292802:00011:00001",
  "USGS:310931081291002:00011:00011",
  "USGS:310931081291002:00011:00001",
  "USGS:311022081304601:00011:00001",
  "USGS:311022081304602:00011:00002",
  "USGS:311022081304602:00011:00001",
  "USGS:311028081285902:00011:00002",
  "USGS:311028081285902:00011:00001",
  "USGS:311051081295501:00011:00001",
  "USGS:311802084192301:00011:00001",
  "USGS:312127084065801:00011:00001",
  "USGS:312232084391701:00011:00001",
  "USGS:312617084110701:00011:00001",
  "USGS:312919084153801:00011:00001",
  "USGS:313118083325401:00011:00002",
  "USGS:313118083325401:00011:00001",
  "USGS:313118083325401:00011:00007",
  "USGS:313118083325401:00011:00011",
  "USGS:313118083325401:00011:00003",
  "USGS:313118083325401:00011:00005",
  "USGS:313118083325401:00011:00004",
  "USGS:313118083325401:00011:00006",
  "USGS:313118083325401:00011:00008",
  "USGS:313118083325401:00011:00009",
  "USGS:313118083325401:00011:00010",
  "USGS:313118083325401:00011:00013",
  "USGS:313118083325401:00011:00014",
  "USGS:313118083325401:00011:00015",
  "USGS:313247084005001:00011:00001",
  "USGS:313808084093601:00011:00001",
  "USGS:320127080511201:00011:00001",
  "USGS:320127080511203:00011:00002",
  "USGS:320127080511203:00011:00001",
  "USGS:320127080511205:00011:00001",
  "USGS:320127080511301:00011:00002",
  "USGS:320127080511301:00011:00001",
  "USGS:320139083511602:00011:00001",
  "USGS:03336645:00011:00002",
  "USGS:03336645:00011:00005",
  "USGS:03336890:00011:00002",
  "USGS:03336890:00011:00001",
  "USGS:03336890:00011:00005",
  "USGS:03336890:00011:00003",
  "USGS:03336900:00011:00002",
  "USGS:03336900:00011:00003",
  "USGS:03336998:00011:00001",
  "USGS:02353265:00011:00002",
  "USGS:02353265:00011:00004",
  "USGS:02353265:00011:00001",
  "USGS:02353400:00011:00003",
  "USGS:02353400:00011:00001",
  "USGS:02353400:00011:00002",
  "USGS:02353500:00011:00005",
  "USGS:02353500:00011:00001",
  "USGS:02353500:00011:00002",
  "USGS:02354350:00011:00005",
  "USGS:02354350:00011:00004",
  "USGS:02354350:00011:00003",
  "USGS:02354475:00011:00002",
  "USGS:02354475:00011:00001",
  "USGS:02354500:00011:00004",
  "USGS:02354500:00011:00001",
  "USGS:02354500:00011:00002",
  "USGS:02354800:00011:00003",
  "USGS:02354800:00011:00002",
  "USGS:02354800:00011:00001",
  "USGS:02355350:00011:00005",
  "USGS:02355350:00011:00002",
  "USGS:02355350:00011:00001",
  "USGS:02355662:00011:00003",
  "USGS:02355662:00011:00002",
  "USGS:02355662:00011:00001",
  "USGS:02356000:00011:00041",
  "USGS:02356000:00011:00006",
  "USGS:02356000:00011:00007",
  "USGS:02356000:00011:00001",
  "USGS:02356000:00011:00002",
  "USGS:02356638:00011:00002",
  "USGS:02356638:00011:00001",
  "USGS:02357000:00011:00008",
  "USGS:02357000:00011:00002",
  "USGS:02357000:00011:00004",
  "USGS:02357000:00011:00007",
  "USGS:02357150:00011:00006",
  "USGS:02357150:00011:00004",
  "USGS:02357150:00011:00002",
  "USGS:02357150:00011:00001",
  "USGS:02379500:00011:00003",
  "USGS:02379500:00011:00001",
  "USGS:02379500:00011:00002",
  "USGS:02380500:00011:00003",
  "USGS:02380500:00011:00001",
  "USGS:02380500:00011:00002",
  "USGS:02381090:00011:00012",
  "USGS:02381090:00011:00002",
  "USGS:02381090:00011:00001",
  "USGS:02381600:00011:00001",
  "USGS:02381600:00011:00002",
  "USGS:02381600:00011:00003",
  "USGS:02382200:00011:00003",
  "USGS:02382200:00011:00001",
  "USGS:02382200:00011:00002",
  "USGS:02382400:00011:00001",
  "USGS:02382500:00011:00021",
  "USGS:02382500:00011:00002",
  "USGS:02382500:00011:00003",
  "USGS:02383500:00011:00010",
  "USGS:02383500:00011:00002",
  "USGS:02383500:00011:00003",
  "USGS:02383520:00011:00001",
  "USGS:02384500:00011:00005",
  "USGS:02384500:00011:00001",
  "USGS:02384500:00011:00002",
  "USGS:02384540:00011:00002",
  "USGS:02384540:00011:00006",
  "USGS:02385170:00011:00003",
  "USGS:02385170:00011:00002",
  "USGS:02385170:00011:00001",
  "USGS:02385500:00011:00003",
  "USGS:02385500:00011:00001",
  "USGS:02385500:00011:00002",
  "USGS:02385800:00011:00005",
  "USGS:02385800:00011:00003",
  "USGS:02385800:00011:00001",
  "USGS:02385800:00011:00002",
  "USGS:02387000:00011:00002",
  "USGS:02387000:00011:00008",
  "USGS:02387010:00011:00001",
  "USGS:02387500:00011:00007",
  "USGS:02387500:00011:00002",
  "USGS:02387500:00011:00003",
  "USGS:02387520:00011:00002",
  "USGS:02387520:00011:00001",
  "USGS:02387600:00011:00003",
  "USGS:02387600:00011:00002",
  "USGS:02387600:00011:00001",
  "USGS:02388320:00011:00001",
  "USGS:02388320:00011:00002",
  "USGS:02388350:00011:00005",
  "USGS:02388350:00011:00004",
  "USGS:02388350:00011:00003",
  "USGS:02388500:00011:00002",
  "USGS:02388500:00011:00003",
  "USGS:02388525:00011:00002",
  "USGS:02388525:00011:00001",
  "USGS:02388975:00011:00003",
  "USGS:02388975:00011:00002",
  "USGS:02388975:00011:00001",
  "USGS:02389150:00011:00002",
  "USGS:02389150:00011:00004",
  "USGS:02389150:00011:00001",
  "USGS:02390000:00011:00005",
  "USGS:02390000:00011:00001",
  "USGS:02390000:00011:00002",
  "USGS:02390050:00011:00004",
  "USGS:02390050:00011:00002",
  "USGS:02390050:00011:00001",
  "USGS:02390140:00011:00005",
  "USGS:02390140:00011:00002",
  "USGS:02390140:00011:00001",
  "USGS:02390475:00011:00003",
  "USGS:02390475:00011:00002",
  "USGS:02390475:00011:00001",
  "USGS:02391540:00011:00005",
  "USGS:02391540:00011:00004",
  "USGS:02391540:00011:00003",
  "USGS:02391840:00011:00003",
  "USGS:02391840:00011:00002",
  "USGS:02391840:00011:00001",
  "USGS:02391860:00011:00003",
  "USGS:02391860:00011:00002",
  "USGS:02391860:00011:00001",
  "USGS:02392000:00011:00026",
  "USGS:02392000:00011:00002",
  "USGS:02392000:00011:00003",
  "USGS:02392360:00011:00005",
  "USGS:02392360:00011:00004",
  "USGS:02392360:00011:00003",
  "USGS:02392780:00011:00006",
  "USGS:02392780:00011:00002",
  "USGS:02392780:00011:00001",
  "USGS:02392950:00011:00013",
  "USGS:02392950:00011:00002",
  "USGS:02392950:00011:00001",
  "USGS:02392975:00011:00013",
  "USGS:02392975:00011:00002",
  "USGS:02392975:00011:00001",
  "USGS:16294100:00011:00002",
  "USGS:16294100:00011:00001",
  "USGS:16294900:00011:00001",
  "USGS:16294900:00011:00002",
  "USGS:16296500:00011:00001",
  "USGS:16296500:00011:00002",
  "USGS:16301050:00011:00001",
  "USGS:09383500:00011:00001",
  "USGS:09383500:00011:00002",
  "USGS:09384000:00011:00004",
  "USGS:09384000:00011:00003",
  "USGS:09384600:00011:00003",
  "USGS:09384600:00011:00001",
  "USGS:09384600:00011:00002",
  "USGS:09385700:00011:00001",
  "USGS:09385700:00011:00002",
  "USGS:09386030:00011:00014",
  "USGS:09386030:00011:00004",
  "USGS:09386030:00011:00003",
  "USGS:09386300:00011:00001",
  "USGS:09386300:00011:00002",
  "USGS:09390500:00011:00001",
  "USGS:09390500:00011:00002",
  "USGS:09394500:00011:00003",
  "USGS:09394500:00011:00001",
  "USGS:09394500:00011:00002",
  "USGS:09396100:00011:00016",
  "USGS:09396100:00011:00001",
  "USGS:09396100:00011:00002",
  "USGS:09396100:00011:00018",
  "USGS:09397000:00011:00001",
  "USGS:09397000:00011:00002",
  "USGS:09397300:00011:00003",
  "USGS:09397300:00011:00022",
  "USGS:09397300:00011:00021",
  "USGS:09397500:00011:00003",
  "USGS:09397500:00011:00001",
  "USGS:09397500:00011:00002",
  "USGS:09398300:00011:00003",
  "USGS:09398300:00011:00004",
  "USGS:09398300:00011:00001",
  "USGS:09398300:00011:00002",
  "USGS:09398300:00011:00016",
  "USGS:09399400:00011:00001",
  "USGS:09399400:00011:00002",
  "USGS:09400350:00011:00001",
  "USGS:09400350:00011:00002",
  "USGS:09400568:00011:00016",
  "USGS:09400568:00011:00002",
  "USGS:09400568:00011:00001",
  "USGS:09400815:00011:00007",
  "USGS:09400815:00011:00001",
  "USGS:09400815:00011:00002",
  "USGS:09400815:00011:00010",
  "USGS:09401110:00011:00002",
  "USGS:09401110:00011:00001",
  "USGS:09401260:00011:00008",
  "USGS:09401260:00011:00007",
  "USGS:09401265:00011:00001",
  "USGS:09401265:00011:00002",
  "USGS:09402000:00011:00009",
  "USGS:09402000:00011:00003",
  "USGS:09402300:00011:00001",
  "USGS:09402300:00011:00002",
  "USGS:09402500:00011:00001",
  "USGS:09402500:00011:00002",
  "USGS:09403850:00011:00001",
  "USGS:09403850:00011:00002",
  "USGS:09404104:00011:00004",
  "USGS:09404104:00011:00001",
  "USGS:09404104:00011:00002",
  "USGS:09404107:00011:00001",
  "USGS:09404107:00011:00002",
  "USGS:09404110:00011:00001",
  "USGS:09404110:00011:00002",
  "USGS:09404115:00011:00001",
  "USGS:09404115:00011:00002",
  "USGS:09404200:00011:00001",
  "USGS:09404200:00011:00003",
  "USGS:09404208:00011:00002",
  "USGS:09404208:00011:00001",
  "USGS:09404222:00011:00001",
  "USGS:09404222:00011:00002",
  "USGS:09404222:00011:00010",
  "USGS:321302082243601:00011:00001",
  "USGS:322036084590301:00011:00001",
  "USGS:322652083033001:00011:00001",
  "USGS:331711081573701:00011:00001",
  "USGS:331944082025501:00011:00011",
  "USGS:331944082025501:00011:00001",
  "USGS:332221081584601:00011:00001",
  "USGS:332221081584602:00011:00001",
  "USGS:332528082003301:00011:00001",
  "USGS:335517084164001:00011:00001",
  "USGS:342922084511601:00011:00001",
  "USGS:344314083433201:00011:00001",
  "USGS:345403085160001:00011:00001",
  "USGS:12413500:00011:00002",
  "USGS:12413500:00011:00001",
  "USGS:12413860:00011:00006",
  "USGS:12413860:00011:00001",
  "USGS:12413875:00011:00002",
  "USGS:12413875:00011:00001",
  "USGS:12414500:00011:00001",
  "USGS:12414500:00011:00002",
  "USGS:12414900:00011:00001",
  "USGS:12414900:00011:00002",
  "USGS:12415070:00011:00001",
  "USGS:12415135:00011:00003",
  "USGS:12415135:00011:00004",
  "USGS:12415135:00011:00001",
  "USGS:12415135:00011:00002",
  "USGS:12415500:00011:00001",
  "USGS:12417610:00011:00006",
  "USGS:12417610:00011:00001",
  "USGS:12417650:00011:00002",
  "USGS:12419000:00011:00001",
  "USGS:12419000:00011:00002",
  "USGS:13032500:00011:00001",
  "USGS:13032500:00011:00002",
  "USGS:13032500:00011:00003",
  "USGS:13037500:00011:00004",
  "USGS:13037500:00011:00005",
  "USGS:13038000:00011:00001",
  "USGS:13038000:00011:00002",
  "USGS:02333500:00011:00015",
  "USGS:02333500:00011:00003",
  "USGS:02333500:00011:00001",
  "USGS:02333500:00011:00002",
  "USGS:02334400:00011:00008",
  "USGS:02334400:00011:00009",
  "USGS:02334400:00011:00006",
  "USGS:02334400:00011:00005",
  "USGS:02334400:00011:00004",
  "USGS:02334400:00011:00023",
  "USGS:02334400:00011:00001",
  "USGS:02334400:00011:00019",
  "USGS:02334401:00011:00001",
  "USGS:02334430:00011:00001",
  "USGS:02334430:00011:00002",
  "USGS:02334430:00011:00003",
  "USGS:02334480:00011:00003",
  "USGS:02334480:00011:00004",
  "USGS:02334480:00011:00002",
  "USGS:02334480:00011:00001",
  "USGS:02334480:00011:00005",
  "USGS:02334578:00011:00004",
  "USGS:02334578:00011:00003",
  "USGS:02334578:00011:00002",
  "USGS:02334578:00011:00001",
  "USGS:02334578:00011:00005",
  "USGS:02334620:00011:00003",
  "USGS:02334620:00011:00001",
  "USGS:02334652:00011:00001",
  "USGS:02334652:00011:00003",
  "USGS:02334653:00011:00004",
  "USGS:02334653:00011:00015",
  "USGS:02334653:00011:00003",
  "USGS:02334653:00011:00002",
  "USGS:02334653:00011:00001",
  "USGS:02334885:00011:00005",
  "USGS:02334885:00011:00016",
  "USGS:02334885:00011:00001",
  "USGS:02334885:00011:00002",
  "USGS:02334885:00011:00017",
  "USGS:02335000:00011:00001",
  "USGS:02335000:00011:00007",
  "USGS:02335000:00011:00002",
  "USGS:02335000:00011:00003",
  "USGS:02335000:00011:00008",
  "USGS:02335000:00011:00009",
  "USGS:02335350:00011:00007",
  "USGS:02335350:00011:00003",
  "USGS:02335350:00011:00002",
  "USGS:02335350:00011:00001",
  "USGS:02335350:00011:00008",
  "USGS:02335450:00011:00011",
  "USGS:02335450:00011:00001",
  "USGS:02335450:00011:00002",
  "USGS:02335580:00011:00011",
  "USGS:02335580:00011:00012",
  "USGS:02335580:00011:00001",
  "USGS:02335700:00011:00005",
  "USGS:02335700:00011:00013",
  "USGS:02335700:00011:00001",
  "USGS:02335700:00011:00002",
  "USGS:02335757:00011:00002",
  "USGS:02335757:00011:00001",
  "USGS:02335790:00011:00005",
  "USGS:02335790:00011:00004",
  "USGS:02335790:00011:00003",
  "USGS:02335810:00011:00009",
  "USGS:02335810:00011:00008",
  "USGS:02335810:00011:00005",
  "USGS:02335810:00011:00006",
  "USGS:02335810:00011:00004",
  "USGS:02335810:00011:00021",
  "USGS:02335810:00011:00001",
  "USGS:02335815:00011:00014",
  "USGS:02335815:00011:00002",
  "USGS:02335815:00011:00001",
  "USGS:023358685:00011:00003",
  "USGS:023358685:00011:00002",
  "USGS:023358685:00011:00001",
  "USGS:02335870:00011:00005",
  "USGS:02335870:00011:00013",
  "USGS:02335870:00011:00001",
  "USGS:02335870:00011:00002",
  "USGS:02335910:00011:00019",
  "USGS:02335910:00011:00009",
  "USGS:02335910:00011:00008",
  "USGS:02335990:00011:00003",
  "USGS:02335990:00011:00001",
  "USGS:02336000:00011:00001",
  "USGS:02336000:00011:00007",
  "USGS:02336000:00011:00006",
  "USGS:02336000:00011:00019",
  "USGS:02336000:00011:00020",
  "USGS:02336030:00011:00004",
  "USGS:02336030:00011:00003",
  "USGS:02336030:00011:00001",
  "USGS:02336030:00011:00005",
  "USGS:02336120:00011:00004",
  "USGS:02336120:00011:00003",
  "USGS:02336120:00011:00002",
  "USGS:02336120:00011:00001",
  "USGS:02336120:00011:00005",
  "USGS:02336120:00011:00006",
  "USGS:02336120:00011:00007",
  "USGS:02336120:00011:00008",
  "USGS:02336152:00011:00004",
  "USGS:02336152:00011:00002",
  "USGS:02336152:00011:00001",
  "USGS:02336152:00011:00005",
  "USGS:02336152:00011:00008",
  "USGS:02336152:00011:00006",
  "USGS:02336152:00011:00007",
  "USGS:023362095:00011:00014",
  "USGS:023362095:00011:00004",
  "USGS:023362095:00011:00001",
  "USGS:023362095:00011:00015",
  "USGS:023362095:00011:00016",
  "USGS:023362095:00011:00017",
  "USGS:023362095:00011:00018",
  "USGS:02336240:00011:00004",
  "USGS:02336240:00011:00002",
  "USGS:02336240:00011:00001",
  "USGS:02336240:00011:00005",
  "USGS:02336240:00011:00006",
  "USGS:02336240:00011:00007",
  "USGS:02336240:00011:00008",
  "USGS:02336300:00011:00006",
  "USGS:02336300:00011:00013",
  "USGS:02336300:00011:00001",
  "USGS:02336300:00011:00002",
  "USGS:02336300:00011:00007",
  "USGS:02336300:00011:00008",
  "USGS:02336300:00011:00009",
  "USGS:02336300:00011:00010",
  "USGS:02336313:00011:00004",
  "USGS:02336313:00011:00003",
  "USGS:02336313:00011:00001",
  "USGS:02336313:00011:00002",
  "USGS:02336313:00011:00005",
  "USGS:02336313:00011:00006",
  "USGS:02336313:00011:00007",
  "USGS:02336313:00011:00008",
  "USGS:02336340:00011:00005",
  "USGS:02336340:00011:00004",
  "USGS:02336340:00011:00001",
  "USGS:02336340:00011:00006",
  "USGS:02336340:00011:00007",
  "USGS:02336340:00011:00008",
  "USGS:02336340:00011:00009",
  "USGS:02336360:00011:00004",
  "USGS:02336360:00011:00003",
  "USGS:02336360:00011:00002",
  "USGS:02336360:00011:00001",
  "USGS:02336360:00011:00005",
  "USGS:02336360:00011:00006",
  "USGS:02336360:00011:00007",
  "USGS:02336360:00011:00008",
  "USGS:02336410:00011:00003",
  "USGS:02336410:00011:00002",
  "USGS:02336410:00011:00001",
  "USGS:02336410:00011:00005",
  "USGS:02336410:00011:00006",
  "USGS:02336410:00011:00007",
  "USGS:02336410:00011:00008",
  "USGS:02336490:00011:00002",
  "USGS:02336490:00011:00003",
  "USGS:02336526:00011:00004",
  "USGS:02336526:00011:00003",
  "USGS:02336526:00011:00002",
  "USGS:02336526:00011:00001",
  "USGS:02336526:00011:00005",
  "USGS:02336526:00011:00006",
  "USGS:02336526:00011:00007",
  "USGS:02336526:00011:00008",
  "USGS:02336635:00011:00015",
  "USGS:02336635:00011:00002",
  "USGS:02336635:00011:00004",
  "USGS:02336728:00011:00003",
  "USGS:02336728:00011:00006",
  "USGS:02336728:00011:00002",
  "USGS:02336728:00011:00001",
  "USGS:02336728:00011:00007",
  "USGS:02336728:00011:00008",
  "USGS:02336728:00011:00009",
  "USGS:02336728:00011:00010",
  "USGS:02336840:00011:00003",
  "USGS:02336840:00011:00002",
  "USGS:02336840:00011:00001",
  "USGS:02336870:00011:00003",
  "USGS:02336870:00011:00002",
  "USGS:02336870:00011:00001",
  "USGS:02336910:00011:00003",
  "USGS:02336910:00011:00002",
  "USGS:02336910:00011:00001",
  "USGS:02336968:00011:00013",
  "USGS:02336968:00011:00002",
  "USGS:02336968:00011:00001",
  "USGS:02336986:00011:00003",
  "USGS:02336986:00011:00002",
  "USGS:02336986:00011:00001",
  "USGS:02337000:00011:00022",
  "USGS:02337000:00011:00008",
  "USGS:02337000:00011:00001",
  "USGS:02337000:00011:00002",
  "USGS:02337040:00011:00003",
  "USGS:02337040:00011:00002",
  "USGS:02337040:00011:00001",
  "USGS:02337170:00011:00010",
  "USGS:02337170:00011:00023",
  "USGS:02337170:00011:00002",
  "USGS:02337170:00011:00003",
  "USGS:02337170:00011:00011",
  "USGS:02337170:00011:00012",
  "USGS:02337170:00011:00013",
  "USGS:02337410:00011:00005",
  "USGS:02337410:00011:00003",
  "USGS:02337410:00011:00002",
  "USGS:02337410:00011:00001",
  "USGS:02337410:00011:00006",
  "USGS:02337410:00011:00007",
  "USGS:02337498:00011:00014",
  "USGS:02337498:00011:00003",
  "USGS:02337498:00011:00002",
  "USGS:02337498:00011:00001",
  "USGS:02337500:00011:00031",
  "USGS:02337500:00011:00001",
  "USGS:02337500:00011:00002",
  "USGS:02338000:00011:00007",
  "USGS:02338000:00011:00002",
  "USGS:02338000:00011:00003",
  "USGS:03274650:00011:00001",
  "USGS:03274650:00011:00002",
  "USGS:03275000:00011:00004",
  "USGS:09404343:00011:00002",
  "USGS:09404343:00011:00001",
  "USGS:09413700:00011:00002",
  "USGS:09413700:00011:00001",
  "USGS:09414900:00011:00002",
  "USGS:09414900:00011:00001",
  "USGS:09415000:00011:00001",
  "USGS:09415000:00011:00002",
  "USGS:09415060:00011:00001",
  "USGS:09415060:00011:00002",
  "USGS:09422500:00011:00001",
  "USGS:09422500:00011:00002",
  "USGS:09423550:00011:00019",
  "USGS:09423550:00011:00001",
  "USGS:09423550:00011:00003",
  "USGS:09423560:00011:00003",
  "USGS:09423560:00011:00001",
  "USGS:09423560:00011:00002",
  "USGS:09424447:00011:00015",
  "USGS:09424447:00011:00001",
  "USGS:09424447:00011:00003",
  "USGS:09424450:00011:00012",
  "USGS:09424450:00011:00001",
  "USGS:09424450:00011:00002",
  "USGS:09424900:00011:00015",
  "USGS:09424900:00011:00013",
  "USGS:09424900:00011:00002",
  "USGS:09424900:00011:00003",
  "USGS:09426000:00011:00016",
  "USGS:09513860:00011:00004",
  "USGS:09426000:00011:00005",
  "USGS:09426620:00011:00001",
  "USGS:09426620:00011:00003",
  "USGS:09428500:00011:00001",
  "USGS:09428500:00011:00004",
  "USGS:09428500:00011:00014",
  "USGS:09428500:00011:00019",
  "USGS:09428505:00011:00001",
  "USGS:09428505:00011:00002",
  "USGS:09428510:00011:00003",
  "USGS:09428510:00011:00001",
  "USGS:09428510:00011:00004",
  "USGS:09429030:00011:00001",
  "USGS:09429030:00011:00002",
  "USGS:09429070:00011:00005",
  "USGS:09429070:00011:00003",
  "USGS:09429070:00011:00001",
  "USGS:09429070:00011:00002",
  "USGS:09439000:00011:00001",
  "USGS:09439000:00011:00002",
  "USGS:09439000:00011:00013",
  "USGS:09442000:00011:00001",
  "USGS:09442000:00011:00002",
  "USGS:09442000:00011:00004",
  "USGS:09442000:00011:00005",
  "USGS:09444200:00011:00003",
  "USGS:09444200:00011:00001",
  "USGS:09444200:00011:00002",
  "USGS:09444500:00011:00001",
  "USGS:09444500:00011:00017",
  "USGS:09447000:00011:00003",
  "USGS:09447000:00011:00001",
  "USGS:09447000:00011:00002",
  "USGS:09447800:00011:00003",
  "USGS:09447800:00011:00001",
  "USGS:09447800:00011:00002",
  "USGS:09448500:00011:00001",
  "USGS:09448500:00011:00021",
  "USGS:09460150:00011:00002",
  "USGS:09460150:00011:00003",
  "USGS:09466500:00011:00001",
  "USGS:09466500:00011:00002",
  "USGS:09468500:00011:00001",
  "USGS:09469000:00011:00003",
  "USGS:09469000:00011:00005",
  "USGS:09469500:00011:00016",
  "USGS:09469500:00011:00001",
  "USGS:09469500:00011:00002",
  "USGS:09470380:00011:00004",
  "USGS:09470380:00011:00002",
  "USGS:09470500:00011:00001",
  "USGS:09470500:00011:00002",
  "USGS:09470700:00011:00012",
  "USGS:09470700:00011:00001",
  "USGS:09470700:00011:00002",
  "USGS:09470750:00011:00012",
  "USGS:09470750:00011:00001",
  "USGS:09470750:00011:00002",
  "USGS:09470800:00011:00004",
  "USGS:09470800:00011:00003",
  "USGS:09470920:00011:00002",
  "USGS:09470920:00011:00012",
  "USGS:09470920:00011:00013",
  "USGS:09470920:00011:00015",
  "USGS:09470920:00011:00016",
  "USGS:09471000:00011:00023",
  "USGS:09471000:00011:00011",
  "USGS:09471000:00011:00008",
  "USGS:09471000:00011:00010",
  "USGS:09471310:00011:00012",
  "USGS:09471310:00011:00001",
  "USGS:09471310:00011:00002",
  "USGS:09471380:00011:00012",
  "USGS:09471380:00011:00001",
  "USGS:09471380:00011:00002",
  "USGS:09471400:00011:00012",
  "USGS:09471400:00011:00001",
  "USGS:09471400:00011:00002",
  "USGS:09471550:00011:00001",
  "USGS:09471550:00011:00002",
  "USGS:09472050:00011:00001",
  "USGS:09472050:00011:00002",
  "USGS:09473000:00011:00003",
  "USGS:09473000:00011:00001",
  "USGS:09473000:00011:00002",
  "USGS:09474000:00011:00022",
  "USGS:09474000:00011:00001",
  "USGS:09474000:00011:00002",
  "USGS:09474000:00011:00010",
  "USGS:09513860:00011:00003",
  "USGS:09475500:00011:00004",
  "USGS:09475500:00011:00003",
  "USGS:09475500:00011:00016",
  "USGS:09478500:00011:00014",
  "USGS:09478500:00011:00017",
  "USGS:09478500:00011:00015",
  "USGS:09479350:00011:00002",
  "USGS:09479350:00011:00001",
  "USGS:09480500:00011:00001",
  "USGS:09480500:00011:00002",
  "USGS:09481000:00011:00001",
  "USGS:09481000:00011:00002",
  "USGS:09481000:00011:00003",
  "USGS:09481740:00011:00001",
  "USGS:09481740:00011:00002",
  "USGS:13075000:00011:00001",
  "USGS:13075000:00011:00002",
  "USGS:13075500:00011:00001",
  "USGS:13075500:00011:00002",
  "USGS:13075910:00011:00001",
  "USGS:13075910:00011:00002",
  "USGS:13075983:00011:00001",
  "USGS:13075983:00011:00002",
  "USGS:13077000:00011:00002",
  "USGS:13077000:00011:00003",
  "USGS:13078000:00011:00001",
  "USGS:13078000:00011:00002",
  "USGS:13081500:00011:00002",
  "USGS:13081500:00011:00003",
  "USGS:13082500:00011:00001",
  "USGS:09509501:00011:00004",
  "USGS:09509502:00011:00001",
  "USGS:09509502:00011:00003",
  "USGS:09510000:00011:00011",
  "USGS:09510000:00011:00010",
  "USGS:09510200:00011:00003",
  "USGS:09510200:00011:00001",
  "USGS:09510200:00011:00002",
  "USGS:09511300:00011:00015",
  "USGS:09511300:00011:00001",
  "USGS:09511300:00011:00016",
  "USGS:09512162:00011:00004",
  "USGS:09512162:00011:00003",
  "USGS:09512165:00011:00002",
  "USGS:09512165:00011:00001",
  "USGS:09512280:00011:00003",
  "USGS:09512280:00011:00001",
  "USGS:09512280:00011:00002",
  "USGS:09512450:00011:00014",
  "USGS:09512450:00011:00001",
  "USGS:09512450:00011:00002",
  "USGS:09512500:00011:00003",
  "USGS:09512500:00011:00001",
  "USGS:09512500:00011:00002",
  "USGS:09512800:00011:00003",
  "USGS:09512800:00011:00001",
  "USGS:09512800:00011:00002",
  "USGS:09513780:00011:00004",
  "USGS:09513780:00011:00002",
  "USGS:09513780:00011:00003",
  "USGS:09514100:00011:00002",
  "USGS:09514100:00011:00001",
  "USGS:09516500:00011:00014",
  "USGS:09516500:00011:00004",
  "USGS:09516500:00011:00003",
  "USGS:09517000:00011:00001",
  "USGS:09517000:00011:00002",
  "USGS:09517000:00011:00021",
  "USGS:09517490:00011:00001",
  "USGS:09517490:00011:00002",
  "USGS:09518500:00011:00004",
  "USGS:09518500:00011:00003",
  "USGS:09519000:00011:00004",
  "USGS:09519000:00011:00003",
  "USGS:09519000:00011:00011",
  "USGS:09519501:00011:00005",
  "USGS:09519501:00011:00004",
  "USGS:09519800:00011:00001",
  "USGS:09519800:00011:00006",
  "USGS:09520280:00011:00014",
  "USGS:09520280:00011:00001",
  "USGS:09520280:00011:00003",
  "USGS:09520500:00011:00001",
  "USGS:09520500:00011:00005",
  "USGS:09522400:00011:00001",
  "USGS:09522400:00011:00002",
  "USGS:09522400:00011:00003",
  "USGS:09522500:00011:00002",
  "USGS:09522500:00011:00006",
  "USGS:09522600:00011:00001",
  "USGS:09522600:00011:00005",
  "USGS:09522650:00011:00001",
  "USGS:09522650:00011:00004",
  "USGS:09522660:00011:00001",
  "USGS:09522660:00011:00002",
  "USGS:09522680:00011:00001",
  "USGS:09522680:00011:00014",
  "USGS:09522680:00011:00002",
  "USGS:09522700:00011:00001",
  "USGS:09522700:00011:00002",
  "USGS:09522700:00011:00022",
  "USGS:09522710:00011:00001",
  "USGS:09522720:00011:00001",
  "USGS:09522730:00011:00001",
  "USGS:09522740:00011:00002",
  "USGS:09522750:00011:00001",
  "USGS:09522760:00011:00001",
  "USGS:09522770:00011:00001",
  "USGS:09522800:00011:00012",
  "USGS:09522800:00011:00001",
  "USGS:09522800:00011:00002",
  "USGS:09522850:00011:00012",
  "USGS:09522850:00011:00013",
  "USGS:09522850:00011:00002",
  "USGS:09522860:00011:00001",
  "USGS:09522880:00011:00001",
  "USGS:09522880:00011:00002",
  "USGS:09522900:00011:00012",
  "USGS:09522900:00011:00001",
  "USGS:09522900:00011:00002",
  "USGS:09525500:00011:00021",
  "USGS:09525500:00011:00002",
  "USGS:09525500:00011:00022",
  "USGS:09526000:00011:00001",
  "USGS:09528200:00011:00002",
  "USGS:09528200:00011:00001",
  "USGS:131610556:00011:00001",
  "USGS:13168500:00011:00014",
  "USGS:13168500:00011:00001",
  "USGS:13168500:00011:00002",
  "USGS:13171500:00011:00001",
  "USGS:13176400:00011:00003",
  "USGS:13176400:00011:00002",
  "USGS:13176400:00011:00001",
  "USGS:13185000:00011:00002",
  "USGS:13185000:00011:00003",
  "USGS:13186000:00011:00002",
  "USGS:13186000:00011:00003",
  "USGS:13190500:00011:00002",
  "USGS:13190500:00011:00003",
  "USGS:13192200:00011:00001",
  "USGS:13192200:00011:00003",
  "USGS:13192200:00011:00002",
  "USGS:13200000:00011:00002",
  "USGS:13200000:00011:00003",
  "USGS:13201500:00011:00004",
  "USGS:13204640:00011:00002",
  "USGS:13204640:00011:00001",
  "USGS:13206000:00011:00001",
  "USGS:13206000:00011:00002",
  "USGS:03337000:00011:00028",
  "USGS:03337000:00011:00001",
  "USGS:03337000:00011:00005",
  "USGS:03337100:00011:00002",
  "USGS:03337100:00011:00001",
  "USGS:03337570:00011:00002",
  "USGS:03337570:00011:00001",
  "USGS:03338780:00011:00003",
  "USGS:03338780:00011:00002",
  "USGS:03339000:00011:00017",
  "USGS:03339000:00011:00005",
  "USGS:03339000:00011:00002",
  "USGS:03339000:00011:00018",
  "USGS:03339000:00011:00019",
  "USGS:03339000:00011:00024",
  "USGS:03339000:00011:00021",
  "USGS:03339000:00011:00032",
  "USGS:03339000:00011:00015",
  "USGS:03339000:00011:00029",
  "USGS:03339000:00011:00030",
  "USGS:03343400:00011:00004",
  "USGS:03343400:00011:00003",
  "USGS:03343805:00011:00003",
  "USGS:03343805:00011:00001",
  "USGS:03343805:00011:00004",
  "USGS:03343805:00011:00005",
  "USGS:03343805:00011:00006",
  "USGS:03343820:00011:00003",
  "USGS:03343820:00011:00001",
  "USGS:03343820:00011:00004",
  "USGS:03345500:00011:00004",
  "USGS:03345500:00011:00002",
  "USGS:03346000:00011:00001",
  "USGS:03346000:00011:00003",
  "USGS:03346500:00011:00001",
  "USGS:03346500:00011:00002",
  "USGS:16019000:00011:00001",
  "USGS:16019000:00011:00002",
  "USGS:16060000:00011:00001",
  "USGS:16060000:00011:00002",
  "USGS:16068000:00011:00001",
  "USGS:16068000:00011:00002",
  "USGS:16071500:00011:00001",
  "USGS:16071500:00011:00002",
  "USGS:16094150:00011:00001",
  "USGS:16097500:00011:00001",
  "USGS:16097500:00011:00002",
  "USGS:16103000:00011:00001",
  "USGS:16103000:00011:00002",
  "USGS:16108000:00011:00002",
  "USGS:16108000:00011:00003",
  "USGS:16200000:00011:00001",
  "USGS:16200000:00011:00013",
  "USGS:16200000:00011:00002",
  "USGS:16200000:00011:00012",
  "USGS:16200000:00011:00014",
  "USGS:16200000:00011:00015",
  "USGS:16208000:00011:00001",
  "USGS:16208000:00011:00002",
  "USGS:16208400:00011:00001",
  "USGS:16210000:00011:00001",
  "USGS:16210100:00011:00001",
  "USGS:16210100:00011:00002",
  "USGS:16210200:00011:00001",
  "USGS:16210200:00011:00005",
  "USGS:16210200:00011:00002",
  "USGS:16210200:00011:00015",
  "USGS:16210200:00011:00003",
  "USGS:16210200:00011:00004",
  "USGS:16210500:00011:00005",
  "USGS:16210500:00011:00002",
  "USGS:16210500:00011:00015",
  "USGS:16210500:00011:00003",
  "USGS:16210500:00011:00004",
  "USGS:16211600:00011:00001",
  "USGS:16211600:00011:00002",
  "USGS:16212480:00011:00001",
  "USGS:16212480:00011:00003",
  "USGS:16212480:00011:00002",
  "USGS:16212480:00011:00004",
  "USGS:16212480:00011:00005",
  "USGS:16212490:00011:00005",
  "USGS:16212490:00011:00002",
  "USGS:16212490:00011:00003",
  "USGS:16212490:00011:00004",
  "USGS:16213000:00011:00002",
  "USGS:16213000:00011:00003",
  "USGS:16226200:00011:00001",
  "USGS:16226200:00011:00008",
  "USGS:16226200:00011:00004",
  "USGS:16226200:00011:00006",
  "USGS:16226200:00011:00002",
  "USGS:16226200:00011:00003",
  "USGS:16226400:00011:00002",
  "USGS:16226400:00011:00004",
  "USGS:16226400:00011:00001",
  "USGS:16226400:00011:00005",
  "USGS:16226400:00011:00015",
  "USGS:16226400:00011:00016",
  "USGS:16227500:00011:00003",
  "USGS:16227500:00011:00004",
  "USGS:16229000:00011:00001",
  "USGS:16229000:00011:00002",
  "USGS:16238000:00011:00001",
  "USGS:16238000:00011:00005",
  "USGS:16238000:00011:00002",
  "USGS:16238000:00011:00003",
  "USGS:16238000:00011:00004",
  "USGS:16238500:00011:00001",
  "USGS:16238500:00011:00012",
  "USGS:16238500:00011:00002",
  "USGS:16240500:00011:00001",
  "USGS:16240500:00011:00013",
  "USGS:16240500:00011:00002",
  "USGS:16240500:00011:00014",
  "USGS:16240500:00011:00015",
  "USGS:16241600:00011:00001",
  "USGS:16241600:00011:00002",
  "USGS:16242500:00011:00002",
  "USGS:16242500:00011:00015",
  "USGS:16242500:00011:00001",
  "USGS:16244000:00011:00001",
  "USGS:16244000:00011:00012",
  "USGS:16244000:00011:00002",
  "USGS:16247100:00011:00001",
  "USGS:16247100:00011:00012",
  "USGS:16247100:00011:00002",
  "USGS:16247100:00011:00014",
  "USGS:16247100:00011:00015",
  "USGS:16254000:00011:00001",
  "USGS:16254000:00011:00002",
  "USGS:16264600:00011:00001",
  "USGS:16275000:00011:00001",
  "USGS:16275000:00011:00002",
  "USGS:16283200:00011:00001",
  "USGS:16284200:00011:00001",
  "USGS:16284200:00011:00002",
  "USGS:03323450:00011:00001",
  "USGS:03323500:00011:00008",
  "USGS:03323500:00011:00016",
  "USGS:03323500:00011:00017",
  "USGS:03323500:00011:00018",
  "USGS:03323500:00011:00019",
  "USGS:03323500:00011:00020",
  "USGS:03323500:00011:00021",
  "USGS:03323500:00011:00022",
  "USGS:03323500:00011:00023",
  "USGS:09528800:00011:00001",
  "USGS:09528800:00011:00004",
  "USGS:09529000:00011:00001",
  "USGS:09529000:00011:00005",
  "USGS:09529150:00011:00001",
  "USGS:09529150:00011:00004",
  "USGS:09529250:00011:00001",
  "USGS:09529250:00011:00004",
  "USGS:09529300:00011:00001",
  "USGS:09529300:00011:00015",
  "USGS:09529420:00011:00001",
  "USGS:09530100:00011:00001",
  "USGS:09536345:00011:00004",
  "USGS:09536345:00011:00001",
  "USGS:09536345:00011:00002",
  "USGS:09536345:00011:00011",
  "USGS:09537200:00011:00004",
  "USGS:09537200:00011:00003",
  "USGS:09537500:00011:00012",
  "USGS:09537500:00011:00001",
  "USGS:09537500:00011:00002",
  "USGS:312101110170601:00011:00001",
  "USGS:322900111153000:00011:00001",
  "USGS:332053110455800:00011:00001",
  "USGS:333806109193500:00011:00013",
  "USGS:333806109193500:00011:00001",
  "USGS:333806109193500:00011:00011",
  "USGS:333806109193500:00011:00012",
  "USGS:335146111280800:00011:00001",
  "AZ011:340553110562745:00011:00001",
  "AZ011:340553110562745:00011:00002",
  "AZ011:340639111162945:00011:00001",
  "AZ011:340639111162945:00011:00002",
  "USGS:340642109501701:00011:00001",
  "USGS:341800110570000:00011:00001",
  "USGS:342059111415500:00011:00001",
  "USGS:342300111054300:00011:00001",
  "USGS:342427111222800:00011:00011",
  "USGS:342427111222800:00011:00001",
  "AZ011:342946111342645:00011:00001",
  "AZ011:342946111342645:00011:00002",
  "USGS:343616111310200:00011:00001",
  "USGS:343636111501400:00011:00001",
  "AZ011:344433111242845:00011:00013",
  "AZ011:344433111242845:00011:00001",
  "AZ011:344433111242845:00011:00002",
  "AZ011:344433111242845:00011:00011",
  "AZ011:344433111242845:00011:00012",
  "USGS:345141111361900:00011:00001",
  "USGS:345603110450301:00011:00002",
  "USGS:350002110355501:00011:00002",
  "USGS:350800112040000:00011:00001",
  "USGS:350802111403400:00011:00001",
  "USGS:350959110562303:00011:00002",
  "USGS:351022111061801:00011:00002",
  "USGS:351214111022101:00011:00002",
  "USGS:351848111323301:00011:00001",
  "USGS:351848111323301:00011:00002",
  "USGS:351907111311601:00011:00001",
  "USGS:351919111311601:00011:00001",
  "USGS:351920111305701:00011:00001",
  "USGS:351932111311601:00011:00001",
  "USGS:352025111332401:00011:00001",
  "USGS:352025111332401:00011:00002",
  "USGS:352500112423000:00011:00001",
  "USGS:360055110304001:00011:00013",
  "USGS:361225110240701:00011:00013",
  "USGS:362936109564101:00011:00013",
  "USGS:363143110355001:00011:00013",
  "USGS:363850110100801:00011:00015",
  "USGS:364338110154601:00011:00013",
  "USGS:365236112442501:00011:00001",
  "USGS:365403112452801:00011:00001",
  "USGS:365602112460201:00011:00001",
  "USGS:03329700:00011:00001",
  "USGS:03329700:00011:00002",
  "USGS:03329900:00011:00001",
  "USGS:03330241:00011:00001",
  "USGS:03330241:00011:00002",
  "USGS:03330500:00011:00001",
  "USGS:03330500:00011:00002",
  "USGS:03331010:00011:00001",
  "USGS:03331040:00011:00001",
  "USGS:03331440:00011:00002",
  "USGS:03331500:00011:00001",
  "USGS:09484550:00011:00002",
  "USGS:09484580:00011:00003",
  "USGS:09484580:00011:00001",
  "USGS:09484580:00011:00002",
  "USGS:09484600:00011:00001",
  "USGS:09484600:00011:00002",
  "USGS:09485000:00011:00001",
  "USGS:09485000:00011:00006",
  "USGS:09485450:00011:00003",
  "USGS:09485450:00011:00004",
  "USGS:09485700:00011:00001",
  "USGS:09485700:00011:00002",
  "USGS:09486055:00011:00001",
  "USGS:09486055:00011:00002",
  "USGS:09486350:00011:00001",
  "USGS:09486350:00011:00002",
  "USGS:09486500:00011:00008",
  "USGS:09486500:00011:00007",
  "USGS:09486520:00011:00015",
  "USGS:09486520:00011:00014",
  "USGS:09486590:00011:00001",
  "USGS:09486590:00011:00002",
  "USGS:09486800:00011:00003",
  "USGS:09486800:00011:00004",
  "USGS:09487000:00011:00001",
  "USGS:09487000:00011:00002",
  "USGS:09489000:00011:00004",
  "USGS:09489000:00011:00003",
  "USGS:09489500:00011:00003",
  "USGS:09489500:00011:00001",
  "USGS:09489500:00011:00002",
  "USGS:09490500:00011:00001",
  "USGS:09490500:00011:00002",
  "USGS:09492400:00011:00001",
  "USGS:09492400:00011:00002",
  "USGS:09494000:00011:00003",
  "USGS:09494000:00011:00001",
  "USGS:09494000:00011:00002",
  "USGS:09496500:00011:00003",
  "USGS:09496500:00011:00001",
  "USGS:09496500:00011:00002",
  "USGS:09497500:00011:00003",
  "USGS:09497500:00011:00001",
  "USGS:09497500:00011:00002",
  "USGS:09497500:00011:00004",
  "USGS:09497700:00011:00011",
  "USGS:09497700:00011:00001",
  "USGS:09497700:00011:00013",
  "USGS:09497800:00011:00003",
  "USGS:09497800:00011:00001",
  "USGS:09497800:00011:00002",
  "USGS:09497980:00011:00003",
  "USGS:09497980:00011:00001",
  "USGS:09497980:00011:00002",
  "USGS:09498400:00011:00014",
  "USGS:09498400:00011:00004",
  "USGS:09498400:00011:00003",
  "USGS:09498500:00011:00003",
  "USGS:09498500:00011:00001",
  "USGS:09498500:00011:00002",
  "USGS:094985005:00011:00001",
  "USGS:094985005:00011:00002",
  "USGS:09498501:00011:00001",
  "USGS:09498501:00011:00002",
  "USGS:09498502:00011:00012",
  "USGS:09498502:00011:00001",
  "USGS:09498502:00011:00002",
  "USGS:09498503:00011:00005",
  "USGS:09498503:00011:00003",
  "USGS:09498503:00011:00004",
  "USGS:09499000:00011:00003",
  "USGS:09499000:00011:00001",
  "USGS:09499000:00011:00002",
  "USGS:09502000:00011:00003",
  "USGS:09502000:00011:00001",
  "USGS:09502000:00011:00002",
  "USGS:09502800:00011:00014",
  "USGS:09502800:00011:00003",
  "USGS:09502800:00011:00004",
  "USGS:09502900:00011:00005",
  "USGS:09502900:00011:00006",
  "USGS:09502960:00011:00016",
  "USGS:09502960:00011:00006",
  "USGS:09502960:00011:00005",
  "USGS:09503000:00011:00002",
  "USGS:09503000:00011:00003",
  "USGS:09503300:00011:00014",
  "USGS:09503300:00011:00001",
  "USGS:09503300:00011:00002",
  "USGS:09503700:00011:00003",
  "USGS:09503700:00011:00001",
  "USGS:09503700:00011:00002",
  "USGS:09504000:00011:00003",
  "USGS:09504000:00011:00001",
  "USGS:09504000:00011:00002",
  "USGS:09504420:00011:00003",
  "USGS:09504420:00011:00001",
  "USGS:09504420:00011:00002",
  "USGS:09504500:00011:00005",
  "USGS:09504500:00011:00004",
  "USGS:09505200:00011:00003",
  "USGS:09505200:00011:00001",
  "USGS:09505200:00011:00002",
  "USGS:09505350:00011:00003",
  "USGS:09505350:00011:00001",
  "USGS:09505350:00011:00002",
  "USGS:09505800:00011:00015",
  "USGS:09505800:00011:00001",
  "USGS:09505800:00011:00002",
  "USGS:09506000:00011:00006",
  "USGS:09506000:00011:00004",
  "USGS:09506000:00011:00005",
  "USGS:09507480:00011:00001",
  "USGS:09507480:00011:00002",
  "USGS:294717092250000:00011:00002",
  "USGS:294717092250000:00011:00001",
  "USGS:294717092250000:00011:00003",
  "USGS:294717092250000:00011:00005",
  "USGS:294717092250000:00011:00004",
  "USGS:294717092250000:00011:00006",
  "USGS:03351060:00011:00002",
  "USGS:03351060:00011:00001",
  "USGS:03351071:00011:00001",
  "USGS:03351072:00011:00002",
  "USGS:03351072:00011:00001",
  "USGS:03351201:00011:00016",
  "USGS:03351201:00011:00015",
  "USGS:03351201:00011:00014",
  "USGS:03351201:00011:00017",
  "USGS:03351201:00011:00001",
  "USGS:03351201:00011:00018",
  "USGS:03351203:00011:00011",
  "USGS:03351203:00011:00001",
  "USGS:03351310:00011:00001",
  "USGS:03351310:00011:00002",
  "USGS:03351500:00011:00001",
  "USGS:03351500:00011:00002",
  "USGS:033521504:00011:00002",
  "USGS:033521504:00011:00001",
  "USGS:03352162:00011:00002",
  "USGS:03352162:00011:00001",
  "USGS:03352500:00011:00001",
  "USGS:03352500:00011:00003",
  "USGS:03352690:00011:00001",
  "USGS:03352695:00011:00001",
  "USGS:03352953:00011:00001",
  "USGS:03352953:00011:00002",
  "USGS:03352972:00011:00001",
  "USGS:03352988:00011:00001",
  "USGS:16301050:00011:00002",
  "USGS:16304200:00011:00001",
  "USGS:16304200:00011:00002",
  "USGS:16325000:00011:00002",
  "USGS:16330000:00011:00001",
  "USGS:16330000:00011:00002",
  "USGS:16343100:00011:00001",
  "USGS:16345000:00011:00001",
  "USGS:16345000:00011:00002",
  "USGS:16400000:00011:00001",
  "USGS:16400000:00011:00002",
  "USGS:16414200:00011:00002",
  "USGS:16414200:00011:00001",
  "USGS:16501200:00011:00002",
  "USGS:16501200:00011:00001",
  "USGS:16508000:00011:00001",
  "USGS:16508000:00011:00002",
  "USGS:16518000:00011:00001",
  "USGS:16518000:00011:00002",
  "USGS:16552800:00011:00001",
  "USGS:16552800:00011:00011",
  "USGS:16587000:00011:00001",
  "USGS:16587000:00011:00002",
  "USGS:16604500:00011:00001",
  "USGS:16604500:00011:00002",
  "USGS:16614000:00011:00001",
  "USGS:16614000:00011:00002",
  "USGS:16618000:00011:00012",
  "USGS:16618000:00011:00001",
  "USGS:16618000:00011:00002",
  "USGS:16620000:00011:00001",
  "USGS:16620000:00011:00002",
  "USGS:16704000:00011:00002",
  "USGS:16704000:00011:00003",
  "USGS:16717000:00011:00001",
  "USGS:16717000:00011:00002",
  "USGS:16720000:00011:00001",
  "USGS:16720000:00011:00002",
  "USGS:16725000:00011:00001",
  "USGS:16725000:00011:00002",
  "USGS:16770500:00011:00001",
  "USGS:16770500:00011:00002",
  "USGS:190423155371501:00011:00001",
  "USGS:194117155174801:00011:00002",
  "USGS:194945155534402:00011:00001",
  "USGS:200518155405801:00011:00001",
  "USGS:203721156151601:00011:00001",
  "USGS:205327156351102:00011:00001",
  "USGS:205405156305401:00011:00001",
  "USGS:205437156310501:00011:00001",
  "USGS:205705156312401:00011:00001",
  "USGS:212359157502601:00011:00001",
  "USGS:212428157511201:00011:00002",
  "USGS:212855157504501:00011:00001",
  "USGS:213016158105901:00011:00001",
  "USGS:213133158014201:00011:00001",
  "USGS:213215157552800:00011:00003",
  "USGS:213237157530701:00011:00001",
  "USGS:213259158035101:00011:00001",
  "USGS:213308158035601:00011:00001",
  "USGS:213335157540601:00011:00001",
  "USGS:213608158011101:00011:00011",
  "USGS:213732158010201:00011:00011",
  "USGS:220356159281401:00011:00001",
  "USGS:220427159300201:00011:00001",
  "USGS:220523159341201:00011:00001",
  "USGS:220541159215901:00011:00001",
  "USGS:03361850:00011:00001",
  "USGS:03361850:00011:00002",
  "USGS:03362000:00011:00013",
  "USGS:03362000:00011:00001",
  "USGS:03362000:00011:00002",
  "USGS:03362500:00011:00001",
  "USGS:03362500:00011:00002",
  "USGS:03363000:00011:00013",
  "USGS:03363000:00011:00001",
  "USGS:03363000:00011:00002",
  "USGS:03363220:00011:00001",
  "USGS:03363400:00011:00001",
  "USGS:03363500:00011:00002",
  "USGS:03363500:00011:00003",
  "USGS:03363900:00011:00012",
  "USGS:03363900:00011:00001",
  "USGS:03363900:00011:00002",
  "USGS:03364000:00011:00001",
  "USGS:03364000:00011:00002",
  "USGS:03364042:00011:00002",
  "USGS:13082500:00011:00002",
  "USGS:13083000:00011:00001",
  "USGS:13083000:00011:00002",
  "USGS:13087900:00011:00003",
  "USGS:13087995:00011:00002",
  "USGS:13087995:00011:00001",
  "USGS:13089500:00011:00004",
  "USGS:13089500:00011:00001",
  "USGS:13090500:00011:00001",
  "USGS:13090500:00011:00002",
  "USGS:13092747:00011:00003",
  "USGS:13092747:00011:00002",
  "USGS:13092747:00011:00001",
  "USGS:13094000:00011:00001",
  "USGS:13094000:00011:00002",
  "USGS:13095175:00011:00002",
  "USGS:13095175:00011:00001",
  "USGS:13095500:00011:00001",
  "USGS:13095500:00011:00002",
  "USGS:13106000:00011:00001",
  "USGS:13106000:00011:00002",
  "USGS:13106500:00011:00001",
  "USGS:13106500:00011:00002",
  "USGS:13108150:00011:00001",
  "USGS:13108150:00011:00002",
  "USGS:13112000:00011:00001",
  "USGS:13112000:00011:00002",
  "USGS:13115000:00011:00001",
  "USGS:13115000:00011:00003",
  "USGS:13116500:00011:00001",
  "USGS:13116500:00011:00002",
  "USGS:13118700:00011:00001",
  "USGS:13118700:00011:00002",
  "USGS:13119000:00011:00001",
  "USGS:13119000:00011:00002",
  "USGS:13120000:00011:00001",
  "USGS:13120000:00011:00002",
  "USGS:13120500:00011:00001",
  "USGS:13120500:00011:00002",
  "USGS:13126000:00011:00001",
  "USGS:13126000:00011:00003",
  "USGS:13127000:00011:00001",
  "USGS:13127000:00011:00002",
  "USGS:13132500:00011:00001",
  "USGS:13132500:00011:00002",
  "USGS:13132513:00011:00001",
  "USGS:13132513:00011:00002",
  "USGS:13132520:00011:00001",
  "USGS:13132520:00011:00002",
  "USGS:13132535:00011:00001",
  "USGS:13132535:00011:00002",
  "USGS:13132565:00011:00002",
  "USGS:13132565:00011:00001",
  "USGS:13135500:00011:00017",
  "USGS:13135500:00011:00001",
  "USGS:13135500:00011:00002",
  "USGS:13135520:00011:00013",
  "USGS:13135520:00011:00002",
  "USGS:13135520:00011:00001",
  "USGS:13137000:00011:00013",
  "USGS:13137000:00011:00001",
  "USGS:13137000:00011:00003",
  "USGS:13137500:00011:00016",
  "USGS:13137500:00011:00001",
  "USGS:13137500:00011:00002",
  "USGS:13138000:00011:00013",
  "USGS:13138000:00011:00002",
  "USGS:13138000:00011:00001",
  "USGS:13138650:00011:00001",
  "USGS:13138650:00011:00002",
  "USGS:13139510:00011:00017",
  "USGS:13139510:00011:00001",
  "USGS:13139510:00011:00003",
  "USGS:13140800:00011:00003",
  "USGS:13140800:00011:00002",
  "USGS:13140800:00011:00001",
  "USGS:13141500:00011:00001",
  "USGS:13141500:00011:00002",
  "USGS:13142500:00011:00001",
  "USGS:13142500:00011:00002",
  "USGS:13147900:00011:00001",
  "USGS:13147900:00011:00002",
  "USGS:13148500:00011:00001",
  "USGS:13148500:00011:00002",
  "USGS:13150430:00011:00003",
  "USGS:13150430:00011:00001",
  "USGS:13150430:00011:00002",
  "USGS:13150430:00011:00016",
  "USGS:13152500:00011:00001",
  "USGS:13152500:00011:00002",
  "USGS:13154500:00011:00001",
  "USGS:13154500:00011:00002",
  "USGS:13154500:00011:00003",
  "USGS:13159800:00011:00001",
  "USGS:13159800:00011:00002",
  "USGS:04099750:00011:00001",
  "USGS:04099750:00011:00002",
  "USGS:04099880:00011:00001",
  "USGS:04100180:00011:00001",
  "USGS:04100220:00011:00002",
  "USGS:04100222:00011:00012",
  "USGS:04100222:00011:00001",
  "USGS:04100222:00011:00002",
  "USGS:04100500:00011:00001",
  "USGS:04100500:00011:00002",
  "USGS:04101000:00011:00001",
  "USGS:04101000:00011:00002",
  "USGS:04101370:00011:00002",
  "USGS:04101370:00011:00001",
  "USGS:04177700:00011:00001",
  "USGS:04177720:00011:00003",
  "USGS:04177720:00011:00001",
  "USGS:04177720:00011:00002",
  "USGS:04179520:00011:00001",
  "USGS:04179520:00011:00002",
  "USGS:04180000:00011:00001",
  "USGS:04180000:00011:00002",
  "USGS:04180500:00011:00001",
  "USGS:04180500:00011:00002",
  "USGS:04180500:00011:00013",
  "USGS:03275000:00011:00003",
  "USGS:03275600:00011:00003",
  "USGS:03275600:00011:00004",
  "USGS:03275990:00011:00001",
  "USGS:03276000:00011:00003",
  "USGS:03276000:00011:00002",
  "USGS:03276500:00011:00003",
  "USGS:03276500:00011:00001",
  "USGS:03276500:00011:00002",
  "USGS:03291780:00011:00001",
  "USGS:03291780:00011:00002",
  "USGS:03294000:00011:00001",
  "USGS:03294000:00011:00002",
  "USGS:03302220:00011:00001",
  "USGS:03302220:00011:00002",
  "USGS:03302680:00011:00002",
  "USGS:03302680:00011:00003",
  "USGS:03302800:00011:00001",
  "USGS:03302800:00011:00002",
  "USGS:03302849:00011:00003",
  "USGS:03303000:00011:00001",
  "USGS:03303000:00011:00002",
  "USGS:03303280:00011:00002",
  "USGS:03303280:00011:00001",
  "USGS:03303300:00011:00001",
  "USGS:03303300:00011:00002",
  "USGS:03304300:00011:00002",
  "USGS:03304300:00011:00001",
  "USGS:03322000:00011:00002",
  "USGS:03322000:00011:00001",
  "USGS:03322011:00011:00002",
  "USGS:03322011:00011:00001",
  "USGS:03322900:00011:00005",
  "USGS:03322900:00011:00001",
  "USGS:03322900:00011:00002",
  "USGS:03322985:00011:00001",
  "USGS:03322985:00011:00002",
  "USGS:10039500:00011:00002",
  "USGS:10039500:00011:00005",
  "USGS:10068500:00011:00001",
  "USGS:10068500:00011:00002",
  "USGS:10092700:00011:00016",
  "USGS:10092700:00011:00001",
  "USGS:10092700:00011:00002",
  "USGS:12305000:00011:00001",
  "USGS:12305000:00011:00002",
  "USGS:12305000:00011:00003",
  "USGS:12306500:00011:00001",
  "USGS:12306500:00011:00002",
  "USGS:12308000:00011:00003",
  "USGS:12308000:00011:00002",
  "USGS:12308000:00011:00001",
  "USGS:12308000:00011:00004",
  "USGS:12308500:00011:00004",
  "USGS:12308500:00011:00001",
  "USGS:12308500:00011:00005",
  "USGS:12309500:00011:00003",
  "USGS:12309500:00011:00002",
  "USGS:12310100:00011:00003",
  "USGS:12310100:00011:00002",
  "USGS:12321500:00011:00001",
  "USGS:12321500:00011:00002",
  "USGS:12322000:00011:00010",
  "USGS:12322000:00011:00024",
  "USGS:12322000:00011:00023",
  "USGS:12322000:00011:00004",
  "USGS:12391950:00011:00002",
  "USGS:12391950:00011:00001",
  "USGS:12392155:00011:00002",
  "USGS:12392155:00011:00001",
  "USGS:12392300:00011:00002",
  "USGS:12393000:00011:00004",
  "USGS:12395000:00011:00001",
  "USGS:12395000:00011:00002",
  "USGS:12395500:00011:00001",
  "USGS:12395500:00011:00002",
  "USGS:12411000:00011:00001",
  "USGS:12411000:00011:00002",
  "USGS:12413000:00011:00001",
  "USGS:12413000:00011:00002",
  "USGS:12413125:00011:00002",
  "USGS:12413125:00011:00001",
  "USGS:12413130:00011:00002",
  "USGS:12413130:00011:00001",
  "USGS:12413131:00011:00001",
  "USGS:12413131:00011:00002",
  "USGS:12413210:00011:00002",
  "USGS:12413210:00011:00001",
  "USGS:12413355:00011:00001",
  "USGS:12413355:00011:00002",
  "USGS:12413370:00011:00014",
  "USGS:12413370:00011:00002",
  "USGS:12413370:00011:00003",
  "USGS:12413370:00011:00015",
  "USGS:12413370:00011:00016",
  "USGS:12413445:00011:00017",
  "USGS:12413445:00011:00002",
  "USGS:12413445:00011:00003",
  "USGS:12413445:00011:00018",
  "USGS:12413445:00011:00016",
  "USGS:12413470:00011:00002",
  "USGS:12413470:00011:00001",
  "USGS:220713159361201:00011:00001",
  "USGS:220739159373001:00011:00001",
  "USGS:220927159355001:00011:00001",
  "USGS:03377500:00011:00003",
  "USGS:03377500:00011:00001",
  "USGS:03377500:00011:00002",
  "USGS:03378000:00011:00001",
  "USGS:03378000:00011:00003",
  "USGS:03378635:00011:00001",
  "USGS:03378635:00011:00003",
  "USGS:03379500:00011:00001",
  "USGS:03379500:00011:00003",
  "USGS:03380500:00011:00002",
  "USGS:03380500:00011:00005",
  "USGS:03381495:00011:00002",
  "USGS:03381500:00011:00002",
  "USGS:03381500:00011:00005",
  "USGS:13038500:00011:00015",
  "USGS:13038500:00011:00001",
  "USGS:13038500:00011:00002",
  "USGS:13039000:00011:00001",
  "USGS:13039000:00011:00002",
  "USGS:13039500:00011:00001",
  "USGS:13039500:00011:00002",
  "USGS:13041010:00011:00002",
  "USGS:13041010:00011:00003",
  "USGS:13042500:00011:00001",
  "USGS:13042500:00011:00002",
  "USGS:13046000:00011:00001",
  "USGS:13046000:00011:00002",
  "USGS:13046995:00011:00002",
  "USGS:13046995:00011:00001",
  "USGS:13047500:00011:00002",
  "USGS:13047500:00011:00003",
  "USGS:13047600:00011:00002",
  "USGS:13047600:00011:00001",
  "USGS:13049500:00011:00001",
  "USGS:13049500:00011:00002",
  "USGS:13050500:00011:00001",
  "USGS:13050500:00011:00002",
  "USGS:13052200:00011:00001",
  "USGS:13052200:00011:00002",
  "USGS:13055000:00011:00002",
  "USGS:13055000:00011:00003",
  "USGS:13055250:00011:00001",
  "USGS:13055250:00011:00004",
  "USGS:13055340:00011:00001",
  "USGS:13055340:00011:00002",
  "USGS:13056500:00011:00001",
  "USGS:13056500:00011:00002",
  "USGS:13056500:00011:00003",
  "USGS:13057000:00011:00015",
  "USGS:13057000:00011:00001",
  "USGS:13057000:00011:00002",
  "USGS:13057132:00011:00002",
  "USGS:13057132:00011:00001",
  "USGS:13057155:00011:00002",
  "USGS:13057155:00011:00001",
  "USGS:13057300:00011:00001",
  "USGS:13057300:00011:00002",
  "USGS:13057500:00011:00001",
  "USGS:13057500:00011:00002",
  "USGS:13057940:00011:00001",
  "USGS:13057940:00011:00002",
  "USGS:13058000:00011:00002",
  "USGS:13058000:00011:00003",
  "USGS:13058510:00011:00001",
  "USGS:13058510:00011:00002",
  "USGS:13058520:00011:00001",
  "USGS:13058520:00011:00002",
  "USGS:13058529:00011:00002",
  "USGS:13058529:00011:00001",
  "USGS:13058530:00011:00001",
  "USGS:13058530:00011:00002",
  "USGS:13060000:00011:00001",
  "USGS:13060000:00011:00002",
  "USGS:13062500:00011:00001",
  "USGS:13062500:00011:00002",
  "USGS:13063000:00011:00001",
  "USGS:13066000:00011:00001",
  "USGS:13066000:00011:00002",
  "USGS:13068300:00011:00002",
  "USGS:13068300:00011:00001",
  "USGS:13068495:00011:00001",
  "USGS:13068495:00011:00002",
  "USGS:13068500:00011:00014",
  "USGS:13068500:00011:00001",
  "USGS:13068500:00011:00002",
  "USGS:13069500:00011:00003",
  "USGS:13069500:00011:00001",
  "USGS:13069500:00011:00002",
  "USGS:13073000:00011:00001",
  "USGS:13073000:00011:00002",
  "USGS:05420400:00011:00001",
  "USGS:05435500:00011:00007",
  "USGS:05435500:00011:00018",
  "USGS:05437050:00011:00004",
  "USGS:05437050:00011:00001",
  "USGS:05437500:00011:00007",
  "USGS:05437500:00011:00006",
  "USGS:05437610:00011:00001",
  "USGS:05437641:00011:00001",
  "USGS:05438030:00011:00002",
  "USGS:05438030:00011:00001",
  "USGS:05438170:00011:00002",
  "USGS:05438170:00011:00001",
  "USGS:05438500:00011:00004",
  "USGS:05438500:00011:00003",
  "USGS:13206305:00011:00002",
  "USGS:13206305:00011:00001",
  "USGS:13213000:00011:00026",
  "USGS:13213000:00011:00002",
  "USGS:13213000:00011:00003",
  "USGS:13213000:00011:00020",
  "USGS:13213000:00011:00025",
  "USGS:13213000:00011:00021",
  "USGS:13213000:00011:00023",
  "USGS:13213000:00011:00022",
  "USGS:13213100:00011:00001",
  "USGS:13213100:00011:00002",
  "USGS:13213100:00011:00003",
  "USGS:13213100:00011:00019",
  "USGS:13213100:00011:00025",
  "USGS:13213100:00011:00020",
  "USGS:13213100:00011:00023",
  "USGS:13213100:00011:00022",
  "USGS:13235000:00011:00001",
  "USGS:13235000:00011:00002",
  "USGS:13236500:00011:00001",
  "USGS:13236500:00011:00002",
  "USGS:13237920:00011:00002",
  "USGS:13237920:00011:00001",
  "USGS:13238500:00011:00001",
  "USGS:13239000:00011:00001",
  "USGS:13239000:00011:00002",
  "USGS:13240000:00011:00001",
  "USGS:13240000:00011:00002",
  "USGS:13246000:00011:00002",
  "USGS:13246000:00011:00003",
  "USGS:13247500:00011:00002",
  "USGS:13247500:00011:00003",
  "USGS:13249500:00011:00002",
  "USGS:13249500:00011:00003",
  "USGS:13250000:00011:00001",
  "USGS:13250000:00011:00002",
  "USGS:13251000:00011:00001",
  "USGS:13251000:00011:00002",
  "USGS:13258500:00011:00001",
  "USGS:13258500:00011:00002",
  "USGS:13265500:00011:00001",
  "USGS:13265500:00011:00002",
  "USGS:13266000:00011:00002",
  "USGS:13266000:00011:00003",
  "USGS:13269000:00011:00001",
  "USGS:13269000:00011:00002",
  "USGS:13269000:00011:00003",
  "USGS:13295000:00011:00002",
  "USGS:13295000:00011:00003",
  "USGS:13296000:00011:00001",
  "USGS:13296000:00011:00002",
  "USGS:13296000:00011:00004",
  "USGS:13296500:00011:00001",
  "USGS:13296500:00011:00002",
  "USGS:13297330:00011:00001",
  "USGS:13297330:00011:00002",
  "USGS:13297355:00011:00001",
  "USGS:13297355:00011:00002",
  "USGS:13302005:00011:00001",
  "USGS:13302005:00011:00002",
  "USGS:13302500:00011:00001",
  "USGS:13302500:00011:00002",
  "USGS:13305000:00011:00002",
  "USGS:13305000:00011:00003",
  "USGS:13305310:00011:00002",
  "USGS:13305310:00011:00001",
  "USGS:13306336:00011:00001",
  "USGS:13306336:00011:00002",
  "USGS:13306370:00011:00001",
  "USGS:13306370:00011:00002",
  "USGS:13306385:00011:00002",
  "USGS:13306385:00011:00001",
  "USGS:13307000:00011:00001",
  "USGS:13307000:00011:00002",
  "USGS:13309220:00011:00001",
  "USGS:13309220:00011:00002",
  "USGS:13310199:00011:00002",
  "USGS:13310199:00011:00001",
  "USGS:13310700:00011:00001",
  "USGS:13310700:00011:00002",
  "USGS:13310800:00011:00002",
  "USGS:13310800:00011:00003",
  "USGS:13310800:00011:00001",
  "USGS:13310800:00011:00004",
  "USGS:13310800:00011:00005",
  "USGS:13311000:00011:00012",
  "USGS:13311000:00011:00001",
  "USGS:13311000:00011:00002",
  "USGS:13311000:00011:00013",
  "USGS:13311000:00011:00014",
  "USGS:13311250:00011:00002",
  "USGS:13311250:00011:00003",
  "USGS:13311250:00011:00001",
  "USGS:13311250:00011:00004",
  "USGS:13311250:00011:00005",
  "USGS:13311450:00011:00002",
  "USGS:13311450:00011:00003",
  "USGS:13311450:00011:00001",
  "USGS:13311450:00011:00004",
  "USGS:13311450:00011:00005",
  "USGS:05531500:00011:00004",
  "USGS:05531500:00011:00003",
  "USGS:05532000:00011:00004",
  "USGS:05532000:00011:00003",
  "USGS:05532500:00011:00004",
  "USGS:05532500:00011:00017",
  "USGS:05532600:00011:00001",
  "USGS:05533000:00011:00001",
  "USGS:05533000:00011:00003",
  "USGS:05533400:00011:00012",
  "USGS:05533400:00011:00005",
  "USGS:05533400:00011:00004",
  "USGS:05533600:00011:00002",
  "USGS:05533600:00011:00001",
  "USGS:05534500:00011:00004",
  "USGS:05534500:00011:00003",
  "USGS:05535000:00011:00005",
  "USGS:05535000:00011:00004",
  "USGS:05535070:00011:00004",
  "USGS:05439000:00011:00001",
  "USGS:05439000:00011:00005",
  "USGS:05439500:00011:00004",
  "USGS:05439500:00011:00003",
  "USGS:05440000:00011:00001",
  "USGS:05440000:00011:00019",
  "USGS:05440700:00011:00009",
  "USGS:05440700:00011:00001",
  "USGS:05440700:00011:00004",
  "USGS:05440700:00011:00002",
  "USGS:05442300:00011:00003",
  "USGS:05442300:00011:00002",
  "USGS:05442300:00011:00001",
  "USGS:05443000:00011:00001",
  "USGS:05443500:00011:00007",
  "USGS:05443500:00011:00006",
  "USGS:05444000:00011:00004",
  "USGS:05444000:00011:00003",
  "USGS:05446500:00011:00006",
  "USGS:05446500:00011:00004",
  "USGS:05447500:00011:00008",
  "USGS:05447500:00011:00006",
  "USGS:05448000:00011:00001",
  "USGS:05448000:00011:00003",
  "USGS:05466000:00011:00001",
  "USGS:05466000:00011:00003",
  "USGS:05466500:00011:00004",
  "USGS:05466500:00011:00015",
  "USGS:05467000:00011:00004",
  "USGS:05467000:00011:00015",
  "USGS:03325000:00011:00005",
  "USGS:03323500:00011:00024",
  "USGS:03323500:00011:00025",
  "USGS:03323583:00011:00001",
  "USGS:03323584:00011:00001",
  "USGS:03323587:00011:00003",
  "USGS:03323587:00011:00007",
  "USGS:03323587:00011:00002",
  "USGS:03323587:00011:00001",
  "USGS:03324000:00011:00028",
  "USGS:03324000:00011:00005",
  "USGS:03324000:00011:00004",
  "USGS:03324000:00011:00003",
  "USGS:03324000:00011:00017",
  "USGS:03324000:00011:00018",
  "USGS:03324000:00011:00019",
  "USGS:03324000:00011:00020",
  "USGS:03324000:00011:00021",
  "USGS:03324000:00011:00022",
  "USGS:03324000:00011:00023",
  "USGS:03324000:00011:00024",
  "USGS:03324000:00011:00025",
  "USGS:03324000:00011:00026",
  "USGS:03324300:00011:00003",
  "USGS:03324300:00011:00001",
  "USGS:03324300:00011:00002",
  "USGS:03324450:00011:00001",
  "USGS:03324500:00011:00003",
  "USGS:03324500:00011:00005",
  "USGS:03324500:00011:00002",
  "USGS:03325000:00011:00026",
  "USGS:05469000:00011:00004",
  "USGS:05469000:00011:00017",
  "USGS:05495500:00011:00004",
  "USGS:05495500:00011:00015",
  "USGS:05512500:00011:00001",
  "USGS:05512500:00011:00005",
  "USGS:05520500:00011:00005",
  "USGS:05520500:00011:00019",
  "USGS:05525000:00011:00006",
  "USGS:05525000:00011:00005",
  "USGS:05525500:00011:00001",
  "USGS:05525500:00011:00003",
  "USGS:05526000:00011:00006",
  "USGS:05526000:00011:00005",
  "USGS:05527000:00011:00002",
  "USGS:05527500:00011:00004",
  "USGS:05527500:00011:00005",
  "USGS:05527500:00011:00020",
  "USGS:05527800:00011:00007",
  "USGS:05527800:00011:00004",
  "USGS:05527800:00011:00003",
  "USGS:05527900:00011:00002",
  "USGS:05527900:00011:00001",
  "USGS:05527905:00011:00002",
  "USGS:05527905:00011:00001",
  "USGS:05527910:00011:00002",
  "USGS:05527910:00011:00001",
  "USGS:05527950:00011:00002",
  "USGS:05527950:00011:00001",
  "USGS:05528000:00011:00006",
  "USGS:03325000:00011:00003",
  "USGS:03325000:00011:00004",
  "USGS:03325000:00011:00002",
  "USGS:03325000:00011:00016",
  "USGS:03325000:00011:00017",
  "USGS:03325000:00011:00018",
  "USGS:03325000:00011:00019",
  "USGS:03325000:00011:00020",
  "USGS:03325000:00011:00021",
  "USGS:03325000:00011:00022",
  "USGS:03325000:00011:00023",
  "USGS:03325000:00011:00024",
  "USGS:03325500:00011:00001",
  "USGS:03325500:00011:00002",
  "USGS:03326500:00011:00001",
  "USGS:03326500:00011:00002",
  "USGS:03326950:00011:00001",
  "USGS:03327000:00011:00003",
  "USGS:03327000:00011:00002",
  "USGS:03327500:00011:00003",
  "USGS:03327500:00011:00001",
  "USGS:03327500:00011:00002",
  "USGS:03328000:00011:00001",
  "USGS:03328000:00011:00002",
  "USGS:03328500:00011:00001",
  "USGS:03328500:00011:00002",
  "USGS:03329000:00011:00002",
  "USGS:03329000:00011:00003",
  "USGS:05387320:00011:00001",
  "USGS:05387405:00011:00001",
  "USGS:05387440:00011:00013",
  "USGS:05528000:00011:00004",
  "USGS:05528000:00011:00003",
  "USGS:05528100:00011:00002",
  "USGS:05528100:00011:00001",
  "USGS:05528500:00011:00001",
  "USGS:05528500:00011:00005",
  "USGS:05529000:00011:00004",
  "USGS:05529000:00011:00003",
  "USGS:05529500:00011:00001",
  "USGS:05529500:00011:00003",
  "USGS:05530000:00011:00001",
  "USGS:05530000:00011:00003",
  "USGS:05530750:00011:00001",
  "USGS:05530990:00011:00006",
  "USGS:05530990:00011:00004",
  "USGS:05530990:00011:00003",
  "USGS:05531015:00011:00001",
  "USGS:05531044:00011:00002",
  "USGS:05531044:00011:00001",
  "USGS:05531175:00011:00002",
  "USGS:05531300:00011:00003",
  "USGS:05531300:00011:00002",
  "USGS:05531300:00011:00001",
  "USGS:05531410:00011:00003",
  "USGS:05531410:00011:00002",
  "USGS:05543010:00011:00001",
  "USGS:05543010:00011:00004",
  "USGS:05543010:00011:00005",
  "USGS:05543010:00011:00006",
  "USGS:05543010:00011:00007",
  "USGS:05387440:00011:00002",
  "USGS:05387490:00011:00001",
  "USGS:05387500:00011:00002",
  "USGS:05387500:00011:00005",
  "USGS:05388250:00011:00002",
  "USGS:05388250:00011:00007",
  "USGS:05388310:00011:00001",
  "USGS:073813375:00011:00001",
  "USGS:073813375:00011:00003",
  "USGS:073813375:00011:00017",
  "USGS:073813375:00011:00018",
  "USGS:13313000:00011:00002",
  "USGS:13313000:00011:00003",
  "USGS:13316500:00011:00001",
  "USGS:13316500:00011:00002",
  "USGS:13317000:00011:00001",
  "USGS:13317000:00011:00002",
  "USGS:13317000:00011:00003",
  "USGS:13317660:00011:00012",
  "USGS:13317660:00011:00001",
  "USGS:13317660:00011:00002",
  "USGS:13336500:00011:00002",
  "USGS:13336500:00011:00003",
  "USGS:13337000:00011:00002",
  "USGS:13337000:00011:00003",
  "USGS:13337500:00011:00001",
  "USGS:13337500:00011:00002",
  "USGS:13338500:00011:00001",
  "USGS:13338500:00011:00002",
  "USGS:13340000:00011:00016",
  "USGS:13340000:00011:00001",
  "USGS:13340000:00011:00002",
  "USGS:13340600:00011:00001",
  "USGS:13340600:00011:00002",
  "USGS:13340600:00011:00003",
  "USGS:13341000:00011:00002",
  "USGS:13341000:00011:00001",
  "USGS:13341000:00011:00005",
  "USGS:13341000:00011:00003",
  "USGS:13341000:00011:00006",
  "USGS:13341050:00011:00001",
  "USGS:13341050:00011:00019",
  "USGS:13341050:00011:00018",
  "USGS:13341050:00011:00020",
  "USGS:13341050:00011:00005",
  "USGS:13341050:00011:00002",
  "USGS:13341050:00011:00003",
  "USGS:13341570:00011:00002",
  "USGS:13341570:00011:00001",
  "USGS:13342295:00011:00002",
  "USGS:13342295:00011:00001",
  "USGS:13342340:00011:00002",
  "USGS:13342340:00011:00001",
  "USGS:13342450:00011:00001",
  "USGS:13342450:00011:00002",
  "USGS:13342500:00011:00001",
  "USGS:13342500:00011:00002",
  "USGS:13342500:00011:00003",
  "USGS:13345000:00011:00001",
  "USGS:13345000:00011:00002",
  "USGS:13346800:00011:00001",
  "USGS:13346800:00011:00002",
  "USGS:431920114062401:00011:00002",
  "USGS:432700112470801:00011:00002",
  "USGS:433705116110601:00011:00001",
  "USGS:434307112382601:00011:00001",
  "USGS:475439116503401:00011:00001",
  "USGS:05577500:00011:00001",
  "USGS:05577500:00011:00003",
  "USGS:05578000:00011:00001",
  "USGS:05578000:00011:00002",
  "USGS:05578300:00011:00005",
  "USGS:05578300:00011:00003",
  "USGS:05578300:00011:00001",
  "USGS:05578500:00011:00001",
  "USGS:05578500:00011:00003",
  "USGS:05579500:00011:00001",
  "USGS:05579500:00011:00003",
  "USGS:05579610:00011:00012",
  "USGS:05579610:00011:00002",
  "USGS:05579610:00011:00001",
  "USGS:05579610:00011:00013",
  "USGS:05579610:00011:00011",
  "USGS:05579610:00011:00007",
  "USGS:05579620:00011:00009",
  "USGS:05579620:00011:00002",
  "USGS:05579620:00011:00001",
  "USGS:05579620:00011:00010",
  "USGS:05579620:00011:00008",
  "USGS:03331500:00011:00002",
  "USGS:03331753:00011:00001",
  "USGS:03331753:00011:00002",
  "USGS:03332555:00011:00001",
  "USGS:03332555:00011:00002",
  "USGS:03332605:00011:00012",
  "USGS:03332605:00011:00001",
  "USGS:03332605:00011:00002",
  "USGS:03333050:00011:00005",
  "USGS:03333050:00011:00004",
  "USGS:03333050:00011:00003",
  "USGS:03333080:00011:00001",
  "USGS:03333270:00011:00001",
  "USGS:03333450:00011:00001",
  "USGS:03333450:00011:00002",
  "USGS:03333700:00011:00001",
  "USGS:03333700:00011:00002",
  "USGS:03334000:00011:00001",
  "USGS:03334000:00011:00002",
  "USGS:03334500:00011:00001",
  "USGS:03334500:00011:00002",
  "USGS:03335000:00011:00001",
  "USGS:03335000:00011:00002",
  "USGS:03335500:00011:00001",
  "USGS:03335500:00011:00002",
  "USGS:03335671:00011:00012",
  "USGS:03335671:00011:00001",
  "USGS:03335671:00011:00002",
  "USGS:033356725:00011:00001",
  "USGS:033356725:00011:00002",
  "USGS:03335673:00011:00001",
  "USGS:03335673:00011:00002",
  "USGS:033356786:00011:00001",
  "USGS:033356786:00011:00002",
  "USGS:03336000:00011:00003",
  "USGS:03336000:00011:00004",
  "USGS:03339273:00011:00001",
  "USGS:03339280:00011:00002",
  "USGS:03339280:00011:00001",
  "USGS:03339500:00011:00003",
  "USGS:03339500:00011:00001",
  "USGS:03339500:00011:00002",
  "USGS:03340500:00011:00005",
  "USGS:03340500:00011:00004",
  "USGS:03340500:00011:00003",
  "USGS:03340800:00011:00003",
  "USGS:03340800:00011:00001",
  "USGS:03340800:00011:00002",
  "USGS:03340870:00011:00001",
  "USGS:03340900:00011:00004",
  "USGS:03340900:00011:00002",
  "USGS:03341300:00011:00003",
  "USGS:03341300:00011:00001",
  "USGS:03341300:00011:00002",
  "USGS:03341500:00011:00001",
  "USGS:03341500:00011:00002",
  "USGS:03342000:00011:00001",
  "USGS:03342000:00011:00002",
  "USGS:03342500:00011:00001",
  "USGS:03342500:00011:00002",
  "USGS:03343010:00011:00012",
  "USGS:03343010:00011:00011",
  "USGS:03343010:00011:00001",
  "USGS:03347000:00011:00001",
  "USGS:03347000:00011:00002",
  "USGS:03348000:00011:00003",
  "USGS:03348000:00011:00001",
  "USGS:03348000:00011:00002",
  "USGS:03348130:00011:00001",
  "USGS:03348130:00011:00002",
  "USGS:03349000:00011:00002",
  "USGS:03349000:00011:00003",
  "USGS:03349210:00011:00001",
  "USGS:03349210:00011:00002",
  "USGS:03349510:00011:00017",
  "USGS:03349510:00011:00001",
  "USGS:03349510:00011:00002",
  "USGS:03350655:00011:00001",
  "USGS:03350655:00011:00002",
  "USGS:03350660:00011:00001",
  "USGS:03350660:00011:00002",
  "USGS:03350700:00011:00003",
  "USGS:03350700:00011:00001",
  "USGS:03350700:00011:00002",
  "USGS:03350800:00011:00012",
  "USGS:03350800:00011:00001",
  "USGS:03350800:00011:00002",
  "USGS:03351000:00011:00002",
  "USGS:03351000:00011:00003",
  "USGS:03351005:00011:00001",
  "USGS:03351007:00011:00011",
  "USGS:03351007:00011:00001",
  "USGS:05595240:00011:00005",
  "USGS:05595700:00011:00003",
  "USGS:05595730:00011:00001",
  "USGS:05595730:00011:00003",
  "USGS:05595765:00011:00002",
  "USGS:05595820:00011:00001",
  "USGS:05595820:00011:00003",
  "USGS:05595860:00011:00002",
  "USGS:05597000:00011:00001",
  "USGS:05597000:00011:00003",
  "USGS:05597500:00011:00001",
  "USGS:05597500:00011:00003",
  "USGS:05599490:00011:00005",
  "USGS:05599490:00011:00006",
  "USGS:05599490:00011:00001",
  "USGS:07020500:00011:00005",
  "USGS:07020500:00011:00002",
  "USGS:07022000:00011:00019",
  "USGS:07022000:00011:00005",
  "USGS:07022000:00011:00002",
  "USGS:374453088261701:00011:00001",
  "USCE:374530089194000:00011:00001",
  "USCE:375405089005000:00011:00001",
  "USCE:380215088574200:00011:00001",
  "USCE:380532088092200:00011:00001",
  "USCE:381115088553800:00011:00001",
  "USCE:381139089531700:00011:00001",
  "USCE:381514089022600:00011:00001",
  "USGS:03382100:00011:00002",
  "USGS:03382100:00011:00007",
  "USGS:03382200:00011:00002",
  "USGS:03384450:00011:00002",
  "USGS:03384450:00011:00007",
  "USGS:03384500:00011:00002",
  "USGS:03384500:00011:00001",
  "USGS:03399800:00011:00001",
  "USGS:03399800:00011:00007",
  "USGS:03611500:00011:00002",
  "USGS:03611500:00011:00006",
  "USGS:03612000:00011:00001",
  "USGS:03612000:00011:00003",
  "USGS:03612500:00011:00001",
  "USGS:03612600:00011:00029",
  "USGS:03612600:00011:00024",
  "USGS:03612600:00011:00012",
  "USGS:03612600:00011:00026",
  "USGS:03612600:00011:00001",
  "USGS:03612600:00011:00030",
  "USGS:03612600:00011:00031",
  "USGS:03612600:00011:00028",
  "USGS:03612600:00011:00034",
  "USGS:03612600:00011:00023",
  "USGS:03612600:00011:00027",
  "USGS:04087440:00011:00001",
  "USGS:05414820:00011:00001",
  "USGS:05414820:00011:00003",
  "USGS:05419000:00011:00004",
  "USGS:05419000:00011:00003",
  "USGS:06814000:00011:00004",
  "USGS:06814000:00011:00003",
  "USGS:06820475:00011:00001",
  "USGS:06827000:00011:00006",
  "USGS:06827000:00011:00005",
  "USGS:06845110:00011:00002",
  "USGS:06845110:00011:00001",
  "USGS:06846500:00011:00007",
  "USGS:06846500:00011:00006",
  "USGS:06847900:00011:00004",
  "USGS:06847900:00011:00003",
  "USGS:06848500:00011:00001",
  "USGS:06848500:00011:00002",
  "USGS:06853500:00011:00005",
  "USGS:06853500:00011:00004",
  "USGS:06853800:00011:00004",
  "USGS:06853800:00011:00003",
  "USGS:06854000:00011:00006",
  "USGS:06854500:00011:00002",
  "USGS:06854500:00011:00006",
  "USGS:06855850:00011:00002",
  "USGS:06855850:00011:00001",
  "USGS:06856000:00011:00001",
  "USGS:06856000:00011:00002",
  "USGS:393423086161001:00011:00001",
  "USGS:394426085080601:00011:00012",
  "USGS:394426085080601:00011:00001",
  "USGS:394632086092701:00011:00001",
  "USGS:394952086110901:00011:00001",
  "USGS:400000086023201:00011:00001",
  "USGS:400541085213701:00011:00001",
  "USGS:03357000:00011:00001",
  "USGS:401532085085301:00011:00001",
  "USGS:402851087213501:00011:00002",
  "USGS:402851087213501:00011:00001",
  "USGS:403407086175701:00011:00001",
  "USGS:405829086175801:00011:00001",
  "USGS:405902087141501:00011:00001",
  "USGS:412350086512801:00011:00001",
  "USGS:413026087213601:00011:00001",
  "USGS:413028087303601:00011:00002",
  "USGS:413028087303601:00011:00001",
  "USGS:413028087303601:00011:00005",
  "USGS:413218087151701:00011:00001",
  "USGS:413339087223001:00011:00002",
  "USGS:413339087223001:00011:00001",
  "USGS:413340087285001:00011:00001",
  "USGS:413340087285001:00011:00014",
  "USGS:414318085200601:00011:00001",
  "USGS:401654088212001:00011:00001",
  "USGS:401654088212004:00011:00001",
  "USCE:401734090040700:00011:00001",
  "USGS:401921089282102:00011:00001",
  "USGS:401921089282103:00011:00001",
  "USCE:401949090534600:00011:00001",
  "USGS:401956088453801:00011:00004",
  "USGS:401956088453801:00011:00003",
  "USGS:401956088453801:00011:00002",
  "USGS:401956088453801:00011:00001",
  "USGS:401956088453801:00011:00005",
  "USGS:401956088453801:00011:00006",
  "USGS:05535070:00011:00003",
  "USGS:05535500:00011:00004",
  "USGS:05535500:00011:00003",
  "USGS:05536000:00011:00006",
  "USGS:05536000:00011:00005",
  "USGS:05536101:00011:00004",
  "USGS:05536101:00011:00002",
  "USGS:05536105:00011:00002",
  "USGS:05536105:00011:00001",
  "USGS:05536118:00011:00001",
  "USGS:05536121:00011:00002",
  "USGS:05536123:00011:00035",
  "USGS:05536137:00011:00001",
  "USGS:05536140:00011:00001",
  "USGS:05536162:00011:00002",
  "USGS:05536162:00011:00001",
  "USGS:05536215:00011:00001",
  "USGS:05536215:00011:00003",
  "USGS:05536235:00011:00004",
  "USGS:05536235:00011:00003",
  "USGS:05536255:00011:00004",
  "USGS:05536255:00011:00003",
  "USGS:05536265:00011:00002",
  "USGS:05536265:00011:00001",
  "USGS:05536275:00011:00005",
  "USGS:05536275:00011:00004",
  "USGS:05536290:00011:00007",
  "USGS:05536290:00011:00004",
  "USGS:05536290:00011:00003",
  "USGS:05536340:00011:00004",
  "USGS:05536340:00011:00003",
  "USGS:05536343:00011:00001",
  "USGS:05536500:00011:00004",
  "USGS:05536500:00011:00003",
  "USGS:05536700:00011:00002",
  "USGS:05536700:00011:00001",
  "USGS:05536890:00011:00020",
  "USGS:05536890:00011:00002",
  "USGS:05536890:00011:00005",
  "USGS:05536890:00011:00006",
  "USGS:05536890:00011:00007",
  "USGS:05536890:00011:00047",
  "USGS:05536890:00011:00003",
  "USGS:05536890:00011:00022",
  "USGS:05536890:00011:00001",
  "USGS:05536995:00011:00017",
  "USGS:05536998:00011:00001",
  "USGS:05536998:00011:00002",
  "USGS:05537500:00011:00004",
  "USGS:05537500:00011:00003",
  "USGS:05537980:00011:00002",
  "USGS:05537980:00011:00003",
  "USGS:05537980:00011:00001",
  "USGS:05538360:00011:00001",
  "USGS:05539000:00011:00004",
  "USGS:05539000:00011:00003",
  "USGS:05539670:00011:00001",
  "USGS:05539900:00011:00004",
  "USGS:05539900:00011:00003",
  "USGS:05540060:00011:00005",
  "USGS:05540060:00011:00006",
  "USGS:05540060:00011:00007",
  "USGS:05540095:00011:00004",
  "USGS:05540095:00011:00003",
  "USGS:05540130:00011:00013",
  "USGS:05540130:00011:00004",
  "USGS:05540130:00011:00003",
  "USGS:05540160:00011:00002",
  "USGS:05540160:00011:00001",
  "USGS:05540195:00011:00004",
  "USGS:05540195:00011:00003",
  "USGS:05540250:00011:00006",
  "USGS:05540250:00011:00005",
  "USGS:05540275:00011:00004",
  "USGS:05540275:00011:00001",
  "USGS:05540290:00011:00003",
  "USGS:05540290:00011:00002",
  "USGS:05540290:00011:00001",
  "USGS:05540500:00011:00005",
  "USGS:05540500:00011:00017",
  "USGS:05541710:00011:00003",
  "USGS:05541710:00011:00001",
  "USGS:05542000:00011:00004",
  "USGS:05542000:00011:00015",
  "USGS:415131088143600:00011:00005",
  "USGS:415300088054600:00011:00001",
  "USGS:415318087362701:00011:00004",
  "USGS:415318087362701:00011:00007",
  "USGS:05449500:00011:00006",
  "USGS:03352988:00011:00002",
  "USGS:03353000:00011:00020",
  "USGS:03353000:00011:00001",
  "USGS:03353000:00011:00002",
  "USGS:03353120:00011:00001",
  "USGS:03353120:00011:00002",
  "USGS:033531908:00011:00002",
  "USGS:033531908:00011:00001",
  "USGS:03353200:00011:00013",
  "USGS:03353200:00011:00022",
  "USGS:03353200:00011:00021",
  "USGS:03353200:00011:00020",
  "USGS:03353200:00011:00001",
  "USGS:03353200:00011:00002",
  "USGS:03353200:00011:00014",
  "USGS:03353200:00011:00015",
  "USGS:03353200:00011:00016",
  "USGS:03353200:00011:00032",
  "USGS:03353200:00011:00034",
  "USGS:03353200:00011:00017",
  "USGS:03353200:00011:00031",
  "USGS:03353200:00011:00033",
  "USGS:03353200:00011:00018",
  "USGS:03353240:00011:00001",
  "USGS:03353450:00011:00005",
  "USGS:03353450:00011:00001",
  "USGS:03353451:00011:00002",
  "USGS:03353451:00011:00001",
  "USGS:03353460:00011:00001",
  "USGS:03353460:00011:00002",
  "USGS:03353494:00011:00002",
  "USGS:03353494:00011:00001",
  "USGS:03353500:00011:00001",
  "USGS:03353500:00011:00002",
  "USGS:03353600:00011:00003",
  "USGS:03353600:00011:00001",
  "USGS:03353600:00011:00002",
  "USGS:033536062:00011:00001",
  "USGS:03353611:00011:00003",
  "USGS:03353611:00011:00002",
  "USGS:03353611:00011:00001",
  "USGS:03353620:00011:00001",
  "USGS:03353620:00011:00002",
  "USGS:03353633:00011:00002",
  "USGS:03353633:00011:00001",
  "USGS:03353637:00011:00003",
  "USGS:03353637:00011:00002",
  "USGS:03353800:00011:00001",
  "USGS:03353800:00011:00002",
  "USGS:03353885:00011:00001",
  "USGS:03353885:00011:00002",
  "USGS:03353890:00011:00003",
  "USGS:03353890:00011:00001",
  "USGS:03353890:00011:00002",
  "USGS:03353910:00011:00001",
  "USGS:03353910:00011:00002",
  "USGS:03354000:00011:00004",
  "USGS:03354000:00011:00003",
  "USGS:03354000:00011:00001",
  "USGS:03354000:00011:00002",
  "USGS:03357000:00011:00002",
  "USGS:03357330:00011:00001",
  "USGS:03357330:00011:00002",
  "USGS:03357350:00011:00001",
  "USGS:03357350:00011:00002",
  "USGS:03357500:00011:00005",
  "USGS:03357500:00011:00003",
  "USGS:03358000:00011:00002",
  "USGS:03358000:00011:00003",
  "USGS:03358900:00011:00001",
  "USGS:03359000:00011:00003",
  "USGS:03359000:00011:00002",
  "USGS:03360000:00011:00001",
  "USGS:03360000:00011:00002",
  "USGS:03360500:00011:00001",
  "USGS:03360500:00011:00002",
  "USGS:03360730:00011:00002",
  "USGS:03360730:00011:00001",
  "USGS:03361000:00011:00003",
  "USGS:03361440:00011:00002",
  "USGS:03361500:00011:00001",
  "USGS:03361500:00011:00002",
  "USGS:03361650:00011:00001",
  "USGS:03361650:00011:00002",
  "USGS:03207965:00011:00002",
  "USGS:03207965:00011:00003",
  "USGS:03207995:00011:00002",
  "USGS:03207995:00011:00001",
  "USGS:03208000:00011:00002",
  "USGS:03209300:00011:00003",
  "USGS:04180610:00011:00001",
  "USGS:04181500:00011:00001",
  "USGS:04181500:00011:00002",
  "USGS:04182000:00011:00002",
  "USGS:04182000:00011:00003",
  "USGS:04182755:00011:00003",
  "USGS:04182755:00011:00007",
  "USGS:04182755:00011:00002",
  "USGS:04182755:00011:00001",
  "USGS:04182769:00011:00002",
  "USGS:04182769:00011:00001",
  "USGS:04182808:00011:00001",
  "USGS:04182808:00011:00002",
  "USGS:04182830:00011:00001",
  "USGS:04182867:00011:00001",
  "USGS:04182867:00011:00002",
  "USGS:04182867:00011:00005",
  "USGS:04182867:00011:00003",
  "USGS:04182867:00011:00004",
  "USGS:04182867:00011:00006",
  "USGS:04182900:00011:00011",
  "USGS:04182900:00011:00001",
  "USGS:04182950:00011:00001",
  "USGS:04182950:00011:00002",
  "USGS:04183000:00011:00001",
  "USGS:04183000:00011:00003",
  "USGS:05515500:00011:00025",
  "USGS:05515500:00011:00001",
  "USGS:05515500:00011:00002",
  "USGS:05515500:00011:00026",
  "USGS:05515500:00011:00029",
  "USGS:05515500:00011:00027",
  "USGS:05515500:00011:00028",
  "USGS:05515500:00011:00030",
  "USGS:05516200:00011:00001",
  "USGS:05516500:00011:00002",
  "USGS:05516500:00011:00005",
  "USGS:05516665:00011:00002",
  "USGS:05516665:00011:00014",
  "USGS:05516665:00011:00001",
  "USGS:05516665:00011:00003",
  "USGS:05516665:00011:00004",
  "USGS:05517000:00011:00014",
  "USGS:05517000:00011:00001",
  "USGS:05517000:00011:00002",
  "USGS:05517000:00011:00012",
  "USGS:05517000:00011:00013",
  "USGS:05517010:00011:00002",
  "USGS:05517500:00011:00001",
  "USGS:05517500:00011:00002",
  "USGS:05517530:00011:00001",
  "USGS:05517530:00011:00002",
  "USGS:05518000:00011:00003",
  "USGS:05518000:00011:00006",
  "USGS:05518000:00011:00001",
  "USGS:05522500:00011:00001",
  "USGS:05522500:00011:00002",
  "USGS:05524500:00011:00003",
  "USGS:05524500:00011:00001",
  "USGS:05524500:00011:00002",
  "USGS:03364042:00011:00001",
  "USGS:05536160:00011:00001",
  "USGS:05536165:00011:00001",
  "USGS:05536179:00011:00005",
  "USGS:05536179:00011:00004",
  "USGS:05536179:00011:00003",
  "USGS:05536179:00011:00001",
  "USGS:05536190:00011:00031",
  "USGS:05536190:00011:00033",
  "USGS:05536190:00011:00030",
  "USGS:05536190:00011:00029",
  "USGS:05536190:00011:00035",
  "USGS:05536190:00011:00032",
  "USGS:05536190:00011:00004",
  "USGS:05536190:00011:00001",
  "USGS:05536190:00011:00002",
  "USGS:05536190:00011:00038",
  "USGS:05536195:00011:00017",
  "USGS:05536195:00011:00019",
  "USGS:05536195:00011:00016",
  "USGS:05536195:00011:00015",
  "USGS:05536195:00011:00014",
  "USGS:05536195:00011:00018",
  "USGS:05536195:00011:00001",
  "USGS:05536195:00011:00002",
  "USGS:05536357:00011:00002",
  "USGS:05536357:00011:00001",
  "USGS:05568615:00011:00008",
  "USGS:05593520:00011:00015",
  "USGS:380626087344401:00011:00001",
  "USGS:380758087551001:00011:00001",
  "USGS:382156085382401:00011:00001",
  "USGS:382323086044501:00011:00001",
  "USGS:383247087361001:00011:00002",
  "USGS:391627085534401:00011:00002",
  "USGS:391627085534401:00011:00001",
  "USGS:392820087242601:00011:00001",
  "USGS:05420680:00011:00002",
  "USGS:05420680:00011:00001",
  "USGS:05420850:00011:00001",
  "USGS:05421000:00011:00002",
  "USGS:05421000:00011:00007",
  "USGS:05421682:00011:00003",
  "USGS:05421682:00011:00001",
  "USGS:05421682:00011:00002",
  "USGS:05421740:00011:00002",
  "USGS:05421740:00011:00001",
  "USGS:05421760:00011:00003",
  "USGS:05421760:00011:00001",
  "USGS:05421760:00011:00002",
  "USGS:05421890:00011:00002",
  "USGS:05422000:00011:00001",
  "USGS:05422000:00011:00003",
  "USGS:05422470:00011:00002",
  "USGS:05422470:00011:00018",
  "USGS:05422560:00011:00002",
  "USGS:05422560:00011:00013",
  "USGS:05422600:00011:00002",
  "USGS:05422600:00011:00013",
  "USGS:05448400:00011:00001",
  "USGS:05449500:00011:00002",
  "USGS:03364200:00011:00001",
  "USGS:03364200:00011:00002",
  "USGS:03364340:00011:00001",
  "USGS:03364500:00011:00014",
  "USGS:03364500:00011:00002",
  "USGS:03364500:00011:00003",
  "USGS:03364650:00011:00001",
  "USGS:03364650:00011:00002",
  "USGS:03365500:00011:00003",
  "USGS:03365500:00011:00001",
  "USGS:03365500:00011:00002",
  "USGS:03366500:00011:00001",
  "USGS:03366500:00011:00002",
  "USGS:03368000:00011:00012",
  "USGS:03368000:00011:00001",
  "USGS:03368000:00011:00002",
  "USGS:03369500:00011:00001",
  "USGS:03369500:00011:00002",
  "USGS:03371500:00011:00001",
  "USGS:03371500:00011:00002",
  "USGS:03372400:00011:00002",
  "USGS:03372500:00011:00001",
  "USGS:03372500:00011:00006",
  "USGS:03372500:00011:00004",
  "USGS:03373500:00011:00003",
  "USGS:03373500:00011:00001",
  "USGS:03373500:00011:00002",
  "USGS:03373508:00011:00001",
  "USGS:03373508:00011:00002",
  "USGS:03373560:00011:00002",
  "USGS:03373560:00011:00001",
  "USGS:03373610:00011:00002",
  "USGS:03373610:00011:00001",
  "USGS:03373686:00011:00002",
  "USGS:03373686:00011:00001",
  "USGS:03373695:00011:00002",
  "USGS:03373695:00011:00001",
  "USGS:03373980:00011:00002",
  "USGS:03373980:00011:00004",
  "USGS:03373980:00011:00003",
  "USGS:03374000:00011:00001",
  "USGS:03374000:00011:00002",
  "USGS:03374100:00011:00019",
  "USGS:03374100:00011:00069",
  "USGS:03374100:00011:00031",
  "USGS:03374100:00011:00013",
  "USGS:03374100:00011:00002",
  "USGS:03374100:00011:00003",
  "USGS:03374100:00011:00004",
  "USGS:03374100:00011:00020",
  "USGS:03374100:00011:00036",
  "USGS:03374100:00011:00055",
  "USGS:03374100:00011:00054",
  "USGS:03374498:00011:00003",
  "USGS:03374500:00011:00005",
  "USGS:03374500:00011:00003",
  "USGS:03374500:00011:00002",
  "USGS:03375500:00011:00001",
  "USGS:03375500:00011:00002",
  "USGS:03376300:00011:00001",
  "USGS:03376300:00011:00002",
  "USGS:03376500:00011:00001",
  "USGS:03376500:00011:00002",
  "USGS:03378500:00011:00011",
  "USGS:03378500:00011:00001",
  "USGS:03378550:00011:00001",
  "USGS:03378550:00011:00002",
  "USGS:04092677:00011:00001",
  "USGS:04092677:00011:00003",
  "USGS:04092677:00011:00002",
  "USGS:04092750:00011:00034",
  "USGS:04092750:00011:00038",
  "USGS:04092750:00011:00028",
  "USGS:04092750:00011:00003",
  "USGS:04092750:00011:00008",
  "USGS:04092750:00011:00036",
  "USGS:04092750:00011:00040",
  "USGS:04092750:00011:00035",
  "USGS:04092750:00011:00037",
  "USGS:04093000:00011:00001",
  "USGS:04093000:00011:00002",
  "USGS:04093100:00011:00001",
  "USGS:04093250:00011:00001",
  "USGS:04094000:00011:00001",
  "USGS:04094000:00011:00002",
  "USGS:04094400:00011:00001",
  "USGS:04094400:00011:00002",
  "USGS:04095090:00011:00030",
  "USGS:04095090:00011:00001",
  "USGS:04095090:00011:00003",
  "USGS:04095090:00011:00002",
  "USGS:04095090:00011:00032",
  "USGS:04095090:00011:00036",
  "USGS:04095090:00011:00031",
  "USGS:04095090:00011:00033",
  "USGS:04095095:00011:00002",
  "USGS:04095096:00011:00001",
  "USGS:04095300:00011:00002",
  "USGS:04095300:00011:00003",
  "USGS:04095380:00011:00001",
  "USGS:04095380:00011:00003",
  "USGS:04095380:00011:00002",
  "USGS:04099510:00011:00013",
  "USGS:04099510:00011:00001",
  "USGS:04099510:00011:00002",
  "USGS:05463500:00011:00001",
  "USGS:05463500:00011:00003",
  "USGS:05464000:00011:00001",
  "USGS:05464000:00011:00003",
  "USGS:05464220:00011:00003",
  "USGS:05464220:00011:00015",
  "USGS:05464315:00011:00001",
  "USGS:05464315:00011:00002",
  "USGS:05464420:00011:00014",
  "USGS:05464420:00011:00001",
  "USGS:05464420:00011:00002",
  "USGS:05464420:00011:00015",
  "USGS:05464500:00011:00025",
  "USGS:05464500:00011:00002",
  "USGS:05464500:00011:00005",
  "USGS:05464500:00011:00024",
  "USCE:381711088521700:00011:00001",
  "USCE:381835088591800:00011:00001",
  "USCE:381926089581400:00011:00001",
  "USCE:382130088350500:00011:00001",
  "USCE:382422089522600:00011:00001",
  "USCE:383025089162400:00011:00001",
  "USCE:383211089225400:00011:00001",
  "USCE:383700089211000:00011:00001",
  "USGS:384312090064701:00011:00001",
  "USGS:384312090064703:00011:00001",
  "USCE:384633089295600:00011:00001",
  "USCE:385521089141200:00011:00001",
  "USCE:385738089052000:00011:00001",
  "USNWS:390855089210900:00011:00001",
  "USCE:390937090365500:00011:00001",
  "USCE:391347088503000:00011:00001",
  "USCE:392430088463500:00011:00001",
  "USCE:394211088231100:00011:00001",
  "USCE:394212090384300:00011:00001",
  "USCE:394352088394300:00011:00001",
  "USCE:394432089340200:00011:00001",
  "USGS:394803088215001:00011:00001",
  "USCE:395035089325000:00011:00001",
  "USCE:395600091245600:00011:00001",
  "USCE:400113090261200:00011:00001",
  "USCE:400129090375400:00011:00001",
  "USCE:400603087355000:00011:00001",
  "USGS:400610088122201:00011:00001",
  "USGS:400641088152501:00011:00001",
  "USCE:400727089590600:00011:00001",
  "USGS:401215088432301:00011:00004",
  "USGS:401215088432301:00011:00003",
  "USGS:401215088432301:00011:00002",
  "USGS:401215088432301:00011:00009",
  "USGS:401215088432301:00011:00005",
  "USGS:401215088432301:00011:00006",
  "USGS:05484900:00011:00001",
  "USGS:05484900:00011:00002",
  "USGS:05485500:00011:00002",
  "USGS:05485500:00011:00005",
  "USGS:05485605:00011:00002",
  "USGS:05485605:00011:00001",
  "USGS:05485640:00011:00001",
  "USGS:05485640:00011:00005",
  "USGS:05486000:00011:00001",
  "USGS:05486000:00011:00003",
  "USGS:05486490:00011:00002",
  "USGS:05486490:00011:00006",
  "USGS:05487470:00011:00001",
  "USGS:05487470:00011:00003",
  "USGS:05487520:00011:00017",
  "USGS:05487520:00011:00016",
  "USGS:05487520:00011:00020",
  "USGS:05487520:00011:00021",
  "USGS:05487520:00011:00022",
  "USGS:05487520:00011:00025",
  "USGS:05487520:00011:00002",
  "USGS:05487980:00011:00002",
  "USGS:415318087362701:00011:00003",
  "USGS:415318087362701:00011:00002",
  "USGS:415318087362701:00011:00001",
  "USGS:415318087362701:00011:00005",
  "USCE:415352090091800:00011:00001",
  "USGS:415356087575000:00011:00003",
  "USGS:415356087575000:00011:00010",
  "USGS:415423088081500:00011:00003",
  "USGS:415457088150600:00011:00008",
  "USGS:415713088284701:00011:00002",
  "USGS:415713088284701:00011:00003",
  "USGS:415713088284701:00011:00001",
  "USGS:415737088031100:00011:00002",
  "USGS:415755087525300:00011:00004",
  "USGS:415801088095700:00011:00003",
  "USGS:415817087591901:00011:00002",
  "USGS:420057088001700:00011:00003",
  "USGS:420354088170500:00011:00004",
  "USGS:420453088043200:00011:00001",
  "USGS:420745088025901:00011:00002",
  "USGS:421036088054501:00011:00001",
  "USGS:421056088380801:00011:00002",
  "USGS:421056088380801:00011:00004",
  "USGS:421056088380801:00011:00001",
  "USGS:421120088281801:00011:00001",
  "USGS:421122088222701:00011:00001",
  "USGS:421122088222702:00011:00001",
  "USGS:421132088085901:00011:00001",
  "USCE:421140088595600:00011:00001",
  "USGS:421145088194801:00011:00001",
  "USGS:421145088194802:00011:00001",
  "USGS:421241088101801:00011:00001",
  "USGS:421321088341101:00011:00001",
  "USGS:421341088283701:00011:00001",
  "USGS:421341088283702:00011:00001",
  "USGS:421341088283703:00011:00001",
  "USGS:421533088421801:00011:00002",
  "USGS:421533088421801:00011:00004",
  "USGS:421533088421801:00011:00001",
  "USGS:421547088142301:00011:00001",
  "USGS:421626088311401:00011:00001",
  "USGS:421626088311402:00011:00001",
  "USGS:421653088370901:00011:00001",
  "USGS:421653088370902:00011:00001",
  "USGS:421653088370903:00011:00001",
  "USGS:421747088270701:00011:00007",
  "USGS:421747088270701:00011:00009",
  "USGS:421747088270701:00011:00005",
  "USGS:421747088270701:00011:00004",
  "USGS:421747088270701:00011:00011",
  "USGS:421747088270701:00011:00008",
  "USGS:421747088270701:00011:00001",
  "USCE:421810089371000:00011:00001",
  "USGS:421820088154501:00011:00001",
  "USGS:421820088154502:00011:00001",
  "USGS:421914088125301:00011:00001",
  "USGS:422032088222001:00011:00001",
  "USGS:422120088330901:00011:00001",
  "USGS:422142088303101:00011:00001",
  "USGS:422142088303102:00011:00001",
  "USGS:422142088303103:00011:00001",
  "USGS:422308088195601:00011:00002",
  "USGS:422308088195601:00011:00004",
  "USGS:422308088195601:00011:00001",
  "USGS:422308088195602:00011:00001",
  "USGS:422308088231001:00011:00001",
  "USGS:02489500:00011:00013",
  "USGS:02489500:00011:00002",
  "USGS:02489500:00011:00012",
  "USGS:02489500:00011:00026",
  "USGS:02489800:00011:00001",
  "USGS:02489800:00011:00002",
  "USGS:02489800:00011:00004",
  "USGS:02489800:00011:00005",
  "USGS:02489800:00011:00003",
  "USGS:02490193:00011:00005",
  "USGS:02490200:00011:00003",
  "USGS:02490200:00011:00001",
  "USGS:02490200:00011:00014",
  "USGS:02491500:00011:00005",
  "USGS:02491500:00011:00004",
  "USGS:02491500:00011:00017",
  "USGS:02492000:00011:00008",
  "USGS:02492000:00011:00002",
  "USGS:02492000:00011:00006",
  "USGS:02492000:00011:00021",
  "USGS:02492100:00011:00003",
  "USGS:06862700:00011:00005",
  "USGS:05451080:00011:00004",
  "USGS:05451080:00011:00003",
  "USGS:05451080:00011:00023",
  "USGS:05451080:00011:00024",
  "USGS:05451080:00011:00005",
  "USGS:05451080:00011:00006",
  "USGS:05451080:00011:00007",
  "USGS:05451210:00011:00004",
  "USGS:05451210:00011:00003",
  "USGS:05451210:00011:00014",
  "USGS:05451210:00011:00008",
  "USGS:05451210:00011:00006",
  "USGS:05451210:00011:00031",
  "USGS:05451210:00011:00009",
  "USGS:05451210:00011:00033",
  "USGS:05451210:00011:00034",
  "USGS:05451210:00011:00012",
  "USGS:05451210:00011:00032",
  "USGS:05451210:00011:00027",
  "USGS:05451500:00011:00001",
  "USGS:05451500:00011:00003",
  "USGS:05451700:00011:00001",
  "USGS:05451700:00011:00003",
  "USGS:05451770:00011:00001",
  "USGS:05451770:00011:00002",
  "USGS:05451900:00011:00001",
  "USGS:05451900:00011:00003",
  "USGS:05452000:00011:00001",
  "USGS:05452000:00011:00003",
  "USGS:05452200:00011:00001",
  "USGS:05452200:00011:00003",
  "USGS:05452500:00011:00002",
  "USGS:05453000:00011:00001",
  "USGS:05453000:00011:00003",
  "USGS:05453100:00011:00001",
  "USGS:05453100:00011:00003",
  "USGS:05453200:00011:00001",
  "USGS:05453520:00011:00002",
  "USGS:05453520:00011:00001",
  "USGS:05453600:00011:00002",
  "USGS:05454000:00011:00001",
  "USGS:05454000:00011:00013",
  "USGS:05454090:00011:00003",
  "USGS:05454090:00011:00002",
  "USGS:05454220:00011:00002",
  "USGS:05454220:00011:00016",
  "USGS:05454300:00011:00001",
  "USGS:05454300:00011:00003",
  "USGS:05454500:00011:00002",
  "USGS:05454500:00011:00008",
  "USGS:05455010:00011:00002",
  "USGS:05455100:00011:00027",
  "USGS:05455100:00011:00001",
  "USGS:05455100:00011:00003",
  "USGS:05455100:00011:00026",
  "USGS:05455230:00011:00001",
  "USGS:05455500:00011:00001",
  "USGS:05455500:00011:00003",
  "USGS:05455700:00011:00001",
  "USGS:05455700:00011:00003",
  "USGS:05457505:00011:00003",
  "USGS:05457505:00011:00001",
  "USGS:05457505:00011:00002",
  "USGS:05457700:00011:00001",
  "USGS:05457700:00011:00003",
  "USGS:05458000:00011:00001",
  "USGS:05458000:00011:00017",
  "USGS:05458300:00011:00013",
  "USGS:05458300:00011:00014",
  "USGS:05458300:00011:00017",
  "USGS:05458300:00011:00018",
  "USGS:05458300:00011:00019",
  "USGS:05458300:00011:00002",
  "USGS:05458300:00011:00001",
  "USGS:05458500:00011:00001",
  "USGS:05458500:00011:00016",
  "USGS:05458900:00011:00001",
  "USGS:05458900:00011:00017",
  "USGS:05459490:00011:00001",
  "USGS:05459500:00011:00001",
  "USGS:05459500:00011:00002",
  "USGS:05460000:00011:00001",
  "USGS:05460400:00011:00003",
  "USGS:05460400:00011:00001",
  "USGS:05460400:00011:00002",
  "USGS:05462000:00011:00002",
  "USGS:05462000:00011:00005",
  "USGS:05463000:00011:00001",
  "USGS:05463000:00011:00017",
  "USGS:05463050:00011:00001",
  "USGS:05463050:00011:00005",
  "USGS:05463050:00011:00017",
  "USGS:06867500:00011:00006",
  "USGS:06868100:00011:00006",
  "USGS:06868100:00011:00001",
  "USGS:06868200:00011:00004",
  "USGS:06868200:00011:00003",
  "USGS:06868850:00011:00002",
  "USGS:06868850:00011:00001",
  "USGS:06869500:00011:00001",
  "USGS:06869500:00011:00002",
  "USGS:06869950:00011:00005",
  "USGS:06869950:00011:00004",
  "USGS:06870200:00011:00002",
  "USGS:06871000:00011:00004",
  "USGS:06871000:00011:00003",
  "USGS:06871500:00011:00004",
  "USGS:06871500:00011:00003",
  "USGS:06872500:00011:00001",
  "USGS:06872500:00011:00002",
  "USGS:06873000:00011:00004",
  "USGS:06873000:00011:00003",
  "USGS:06873460:00011:00004",
  "USGS:06873460:00011:00003",
  "USGS:06874000:00011:00015",
  "USGS:06874000:00011:00001",
  "USGS:06874000:00011:00002",
  "USGS:06875900:00011:00004",
  "USGS:06875900:00011:00003",
  "USGS:06876000:00011:00002",
  "USGS:06876000:00011:00006",
  "USGS:05464695:00011:00003",
  "USGS:05464695:00011:00001",
  "USGS:05464695:00011:00002",
  "USGS:05464780:00011:00003",
  "USGS:05464780:00011:00001",
  "USGS:05464780:00011:00002",
  "USGS:05464942:00011:00004",
  "USGS:05464942:00011:00003",
  "USGS:05465000:00011:00001",
  "USGS:05465000:00011:00003",
  "USGS:05465500:00011:00042",
  "USGS:05465500:00011:00002",
  "USGS:05465500:00011:00008",
  "USGS:05465500:00011:00041",
  "USGS:05465500:00011:00023",
  "USGS:05465700:00011:00001",
  "USGS:05465700:00011:00002",
  "USGS:05469860:00011:00001",
  "USGS:05469990:00011:00001",
  "USGS:05470000:00011:00001",
  "USGS:05470000:00011:00002",
  "USGS:05470500:00011:00001",
  "USGS:05470500:00011:00002",
  "USGS:05471000:00011:00001",
  "USGS:05471000:00011:00002",
  "USGS:05471050:00011:00001",
  "USGS:05471050:00011:00010",
  "USGS:05471200:00011:00001",
  "USGS:05471200:00011:00014",
  "USGS:05471500:00011:00001",
  "USGS:05471500:00011:00003",
  "USGS:05472500:00011:00001",
  "USGS:05472500:00011:00003",
  "USGS:05473065:00011:00003",
  "USGS:05473065:00011:00001",
  "USGS:05473065:00011:00002",
  "USGS:05473400:00011:00001",
  "USGS:05473400:00011:00004",
  "USGS:05473450:00011:00002",
  "USGS:05473450:00011:00001",
  "USGS:05474000:00011:00002",
  "USGS:05474000:00011:00008",
  "USGS:05476590:00011:00002",
  "USGS:05476590:00011:00001",
  "USGS:05476590:00011:00015",
  "USGS:05476750:00011:00001",
  "USGS:05476750:00011:00003",
  "USGS:05478265:00011:00012",
  "USGS:05478265:00011:00001",
  "USGS:05478265:00011:00015",
  "USGS:05479000:00011:00001",
  "USGS:05479000:00011:00003",
  "USGS:05480500:00011:00001",
  "USGS:05480500:00011:00003",
  "USGS:05480820:00011:00003",
  "USGS:05480820:00011:00002",
  "USGS:05480820:00011:00001",
  "USGS:05480820:00011:00015",
  "USGS:05481000:00011:00016",
  "USGS:05481000:00011:00001",
  "USGS:05481000:00011:00003",
  "USGS:05481000:00011:00017",
  "USGS:05481300:00011:00001",
  "USGS:05481300:00011:00003",
  "USGS:05481510:00011:00001",
  "USGS:05481650:00011:00002",
  "USGS:05481650:00011:00008",
  "USGS:05481950:00011:00001",
  "USGS:05481950:00011:00003",
  "USGS:05482000:00011:00020",
  "USGS:05482000:00011:00002",
  "USGS:05482000:00011:00017",
  "USGS:05482000:00011:00021",
  "USGS:05482300:00011:00018",
  "USGS:05482300:00011:00001",
  "USGS:05482300:00011:00004",
  "USGS:05482300:00011:00016",
  "USGS:05482315:00011:00003",
  "USGS:05482500:00011:00017",
  "USGS:05482500:00011:00001",
  "USGS:05482500:00011:00003",
  "USGS:05482500:00011:00015",
  "USGS:05483318:00011:00001",
  "USGS:05483349:00011:00003",
  "USGS:05483450:00011:00002",
  "USGS:05483450:00011:00008",
  "USGS:05483470:00011:00005",
  "USGS:05483600:00011:00023",
  "USGS:05483600:00011:00002",
  "USGS:05483600:00011:00008",
  "USGS:05483600:00011:00021",
  "USGS:05484000:00011:00001",
  "USGS:05484000:00011:00003",
  "USGS:05484500:00011:00028",
  "USGS:05484500:00011:00001",
  "USGS:05484500:00011:00003",
  "USGS:05484500:00011:00018",
  "USGS:05484600:00011:00002",
  "USGS:05484600:00011:00001",
  "USGS:05484650:00011:00012",
  "USGS:05484650:00011:00013",
  "USGS:05484800:00011:00001",
  "USGS:05484800:00011:00002",
  "USGS:06891080:00011:00002",
  "USGS:06891080:00011:00001",
  "USGS:06891080:00011:00003",
  "USGS:06891200:00011:00001",
  "USGS:06891260:00011:00002",
  "USGS:06891260:00011:00001",
  "USGS:06891478:00011:00013",
  "USGS:06891478:00011:00001",
  "USGS:06891500:00011:00019",
  "USGS:06891500:00011:00018",
  "USGS:06891500:00011:00001",
  "USGS:06891500:00011:00002",
  "USGS:06891810:00011:00002",
  "USGS:06891810:00011:00001",
  "USGS:06892000:00011:00001",
  "USGS:06892000:00011:00002",
  "USGS:06892350:00011:00018",
  "USGS:06892350:00011:00064",
  "USGS:05579620:00011:00005",
  "USGS:05579624:00011:00001",
  "USGS:05579624:00011:00008",
  "USGS:05579624:00011:00005",
  "USGS:05579624:00011:00002",
  "USGS:05579624:00011:00003",
  "USGS:05579630:00011:00005",
  "USGS:05579630:00011:00002",
  "USGS:05579630:00011:00001",
  "USGS:05579630:00011:00006",
  "USGS:05579630:00011:00008",
  "USGS:05579630:00011:00009",
  "USGS:05579630:00011:00007",
  "USGS:05579630:00011:00022",
  "USGS:05579630:00011:00021",
  "USGS:05579630:00011:00025",
  "USGS:05579630:00011:00016",
  "USGS:05579725:00011:00002",
  "USGS:05579725:00011:00001",
  "USGS:05580000:00011:00004",
  "USGS:05580000:00011:00003",
  "USGS:05580950:00011:00001",
  "USGS:05580950:00011:00003",
  "USGS:05582000:00011:00005",
  "USGS:05582000:00011:00004",
  "USGS:05583000:00011:00005",
  "USGS:05583000:00011:00019",
  "USGS:05584500:00011:00007",
  "USGS:05584500:00011:00004",
  "USGS:05585000:00011:00005",
  "USGS:05585000:00011:00020",
  "USGS:05585500:00011:00032",
  "USGS:05586100:00011:00034",
  "USGS:05586100:00011:00017",
  "USGS:05586300:00011:00020",
  "USGS:05586300:00011:00028",
  "USGS:05586300:00011:00001",
  "USGS:05586300:00011:00021",
  "USGS:05586300:00011:00023",
  "USGS:05586300:00011:00022",
  "USGS:05586300:00011:00024",
  "USGS:05586300:00011:00017",
  "USGS:05586300:00011:00054",
  "USGS:05586300:00011:00058",
  "USGS:05586300:00011:00055",
  "USGS:05586300:00011:00025",
  "USGS:05586300:00011:00016",
  "USGS:05586300:00011:00050",
  "USGS:05586300:00011:00015",
  "USGS:05587000:00011:00004",
  "USGS:05587000:00011:00003",
  "USGS:05587060:00011:00001",
  "USGS:05587450:00011:00016",
  "USGS:05587450:00011:00002",
  "USGS:05587498:00011:00001",
  "USGS:05587900:00011:00001",
  "USGS:05587900:00011:00003",
  "USGS:05588000:00011:00001",
  "USGS:05588000:00011:00003",
  "USGS:05590050:00011:00003",
  "USGS:05590050:00011:00002",
  "USGS:05590050:00011:00001",
  "USGS:05590520:00011:00002",
  "USGS:05590520:00011:00001",
  "USGS:05590800:00011:00001",
  "USGS:05590800:00011:00003",
  "USGS:05590950:00011:00002",
  "USGS:05590950:00011:00001",
  "USGS:05591200:00011:00005",
  "USGS:05591200:00011:00002",
  "USGS:05591550:00011:00004",
  "USGS:05591550:00011:00002",
  "USGS:05591700:00011:00004",
  "USGS:05591700:00011:00002",
  "USGS:05592000:00011:00001",
  "USGS:05592000:00011:00005",
  "USGS:05592050:00011:00004",
  "USGS:05592050:00011:00002",
  "USGS:05592100:00011:00005",
  "USGS:05592100:00011:00002",
  "USGS:05592500:00011:00004",
  "USGS:05592500:00011:00002",
  "USGS:05592575:00011:00001",
  "USGS:05592575:00011:00003",
  "USGS:05592800:00011:00004",
  "USGS:05592800:00011:00002",
  "USGS:05592900:00011:00004",
  "USGS:05592900:00011:00002",
  "USGS:05593000:00011:00005",
  "USGS:05593000:00011:00002",
  "USGS:05593020:00011:00002",
  "USGS:05593575:00011:00001",
  "USGS:05593575:00011:00003",
  "USGS:05593900:00011:00001",
  "USGS:05593900:00011:00003",
  "USGS:05593945:00011:00002",
  "USGS:05593945:00011:00001",
  "USGS:05594000:00011:00004",
  "USGS:05594000:00011:00003",
  "USGS:05594100:00011:00005",
  "USGS:05594100:00011:00002",
  "USGS:05594450:00011:00001",
  "USGS:05594450:00011:00003",
  "USGS:05594800:00011:00001",
  "USGS:05594800:00011:00003",
  "USGS:05595000:00011:00004",
  "USGS:05595000:00011:00001",
  "USGS:05595000:00011:00002",
  "USGS:05595200:00011:00001",
  "USGS:05595200:00011:00003",
  "USGS:07140850:00011:00004",
  "USGS:07140850:00011:00002",
  "USGS:07140880:00011:00001",
  "USGS:07140880:00011:00002",
  "USGS:07140885:00011:00002",
  "USGS:07140885:00011:00001",
  "USGS:07140890:00011:00001",
  "USGS:07140890:00011:00002",
  "USGS:07140900:00011:00001",
  "USGS:07140900:00011:00002",
  "USGS:07141000:00011:00001",
  "USGS:03209300:00011:00002",
  "USGS:03209500:00011:00003",
  "USGS:03209500:00011:00005",
  "USGS:03209500:00011:00002",
  "USGS:03209800:00011:00002",
  "USGS:03210000:00011:00003",
  "USGS:03210000:00011:00006",
  "USGS:03210000:00011:00002",
  "USGS:03211000:00011:00002",
  "USGS:03211000:00011:00001",
  "USGS:03211500:00011:00002",
  "USGS:03212500:00011:00006",
  "USGS:03212500:00011:00002",
  "USGS:05389000:00011:00001",
  "USGS:05389000:00011:00002",
  "USGS:05389400:00011:00002",
  "USGS:05389400:00011:00001",
  "USGS:05389500:00011:00002",
  "USGS:05389500:00011:00004",
  "USGS:05411500:00011:00001",
  "USGS:05411600:00011:00003",
  "USGS:05411600:00011:00001",
  "USGS:05411600:00011:00002",
  "USGS:05411850:00011:00002",
  "USGS:05411850:00011:00001",
  "USGS:05411900:00011:00001",
  "USGS:05411900:00011:00002",
  "USGS:05412020:00011:00001",
  "USGS:05412020:00011:00002",
  "USGS:05412340:00011:00003",
  "USGS:05412340:00011:00001",
  "USGS:05412340:00011:00002",
  "USGS:05412400:00011:00004",
  "USGS:05412400:00011:00003",
  "USGS:05412500:00011:00021",
  "USGS:05412500:00011:00002",
  "USGS:05412500:00011:00007",
  "USGS:05412500:00011:00020",
  "USGS:05414400:00011:00001",
  "USGS:05416900:00011:00002",
  "USGS:05416900:00011:00001",
  "USGS:05418110:00011:00005",
  "USGS:05418110:00011:00003",
  "USGS:05418110:00011:00001",
  "USGS:05418110:00011:00002",
  "USGS:05418110:00011:00007",
  "USGS:05418110:00011:00006",
  "USGS:05418400:00011:00017",
  "USGS:05418400:00011:00021",
  "USGS:05418400:00011:00002",
  "USGS:05418400:00011:00001",
  "USGS:05418400:00011:00022",
  "USGS:05418400:00011:00024",
  "USGS:05418400:00011:00023",
  "USGS:05418400:00011:00025",
  "USGS:05418400:00011:00027",
  "USGS:05418400:00011:00028",
  "USGS:05418400:00011:00026",
  "USGS:05418400:00011:00019",
  "USGS:05418400:00011:00018",
  "USGS:05418400:00011:00029",
  "USGS:05418500:00011:00002",
  "USGS:05418500:00011:00008",
  "USGS:05418720:00011:00013",
  "USGS:05418720:00011:00018",
  "USGS:05418720:00011:00002",
  "USGS:05418720:00011:00015",
  "USGS:05418720:00011:00014",
  "USGS:05418720:00011:00012",
  "USGS:05420460:00011:00019",
  "USGS:05420460:00011:00001",
  "USGS:05420500:00011:00024",
  "USGS:05420500:00011:00002",
  "USGS:05420500:00011:00005",
  "USGS:422308088231002:00011:00001",
  "USGS:422308088264201:00011:00001",
  "USGS:422358088360201:00011:00001",
  "USGS:422433088140601:00011:00001",
  "USGS:422704088385301:00011:00001",
  "USGS:422704088385302:00011:00001",
  "USGS:422803087475301:00011:00001",
  "USGS:422803087475302:00011:00001",
  "USGS:422803087475303:00011:00001",
  "USGS:422803087475304:00011:00001",
  "USGS:422803087475305:00011:00001",
  "USGS:422828088333301:00011:00001",
  "USGS:422834088255800:00011:00001",
  "USGS:422845088285401:00011:00001",
  "USGS:422848088191001:00011:00002",
  "USGS:422848088191001:00011:00004",
  "USGS:422848088191001:00011:00001",
  "USGS:422848088191002:00011:00001",
  "USGS:422848088191003:00011:00001",
  "USGS:422858088235601:00011:00001",
  "USGS:422925088255401:00011:00001",
  "USGS:422925088255402:00011:00001",
  "USGS:55559999:00011:00003",
  "USGS:03611260:00011:00001",
  "USGS:03611260:00011:00003",
  "USGS:07157500:00011:00005",
  "USGS:07157500:00011:00004",
  "USGS:07157740:00011:00010",
  "USGS:07165750:00011:00002",
  "USGS:07165750:00011:00001",
  "USGS:07166500:00011:00001",
  "USGS:07166500:00011:00002",
  "USGS:07167500:00011:00004",
  "USGS:07167500:00011:00003",
  "USGS:07169500:00011:00001",
  "USGS:07169500:00011:00002",
  "USGS:07169800:00011:00001",
  "USGS:07169800:00011:00002",
  "USGS:07170500:00011:00001",
  "USGS:07170500:00011:00002",
  "USGS:07170700:00011:00002",
  "USGS:07170990:00011:00002",
  "USGS:07170990:00011:00001",
  "USGS:07172000:00011:00001",
  "USGS:07172000:00011:00002",
  "USGS:07179300:00011:00002",
  "USGS:05543010:00011:00008",
  "USGS:05543010:00011:00010",
  "USGS:05543010:00011:00009",
  "USGS:05543010:00011:00012",
  "USGS:05543500:00011:00007",
  "USGS:05543500:00011:00004",
  "USGS:05547000:00011:00003",
  "USGS:05547500:00011:00003",
  "USGS:05548000:00011:00003",
  "USGS:05548030:00011:00002",
  "USGS:05548030:00011:00001",
  "USGS:05548105:00011:00003",
  "USGS:05548105:00011:00002",
  "USGS:05548105:00011:00001",
  "USGS:05548280:00011:00007",
  "USGS:05548280:00011:00004",
  "USGS:05548280:00011:00003",
  "USGS:05548500:00011:00003",
  "USGS:05549000:00011:00001",
  "USGS:05549000:00011:00002",
  "USGS:05549500:00011:00003",
  "USGS:05549501:00011:00001",
  "USGS:05550000:00011:00004",
  "USGS:05550000:00011:00003",
  "USGS:05550001:00011:00003",
  "USGS:05550001:00011:00002",
  "USGS:05550300:00011:00003",
  "USGS:05550300:00011:00002",
  "USGS:05550300:00011:00001",
  "USGS:05550500:00011:00004",
  "USGS:05550500:00011:00003",
  "USGS:05551000:00011:00007",
  "USGS:05551000:00011:00006",
  "USGS:05551001:00011:00001",
  "USGS:05551200:00011:00008",
  "USGS:05551200:00011:00004",
  "USGS:05551200:00011:00003",
  "USGS:05551330:00011:00003",
  "USGS:05551330:00011:00002",
  "USGS:05551330:00011:00001",
  "USGS:05551540:00011:00002",
  "USGS:05551540:00011:00001",
  "USGS:05551545:00011:00001",
  "USGS:05551580:00011:00002",
  "USGS:05551580:00011:00001",
  "USGS:05551580:00011:00004",
  "USGS:05551580:00011:00007",
  "USGS:05551580:00011:00006",
  "USGS:05551581:00011:00001",
  "USGS:05551582:00011:00001",
  "USGS:05551675:00011:00003",
  "USGS:05551675:00011:00002",
  "USGS:05551675:00011:00001",
  "USGS:05551700:00011:00004",
  "USGS:05551700:00011:00003",
  "USGS:05552500:00011:00007",
  "USGS:05552500:00011:00004",
  "USGS:05554300:00011:00002",
  "USGS:05554300:00011:00001",
  "USGS:05554300:00011:00006",
  "USGS:05554300:00011:00003",
  "USGS:05554500:00011:00005",
  "USGS:05554500:00011:00004",
  "USGS:05555300:00011:00004",
  "USGS:05555300:00011:00017",
  "USGS:05556500:00011:00001",
  "USGS:05556500:00011:00006",
  "USGS:05558300:00011:00032",
  "USGS:05558300:00011:00029",
  "USGS:05558300:00011:00027",
  "USGS:05558300:00011:00028",
  "USGS:05560500:00011:00001",
  "USGS:05560500:00011:00003",
  "USGS:05561500:00011:00001",
  "USGS:05561500:00011:00003",
  "USGS:05567500:00011:00004",
  "USGS:05567500:00011:00017",
  "USGS:05568000:00011:00001",
  "USGS:05568000:00011:00006",
  "USGS:05568500:00011:00030",
  "USGS:05568500:00011:00006",
  "USGS:05568500:00011:00022",
  "USGS:05568800:00011:00008",
  "USGS:05568800:00011:00007",
  "USGS:05569500:00011:00004",
  "USGS:05569500:00011:00015",
  "USGS:05570000:00011:00004",
  "USGS:05570000:00011:00017",
  "USGS:05570910:00011:00001",
  "USGS:05570910:00011:00003",
  "USGS:05572000:00011:00003",
  "USGS:05572000:00011:00008",
  "USGS:05573540:00011:00004",
  "USGS:05573540:00011:00003",
  "USGS:05575550:00011:00002",
  "USGS:05575550:00011:00001",
  "USGS:05575550:00011:00004",
  "USGS:05575550:00011:00003",
  "USGS:05576000:00011:00004",
  "USGS:05576000:00011:00017",
  "USGS:05576022:00011:00001",
  "USGS:05576250:00011:00002",
  "USGS:05576250:00011:00001",
  "USGS:05576500:00011:00004",
  "USGS:05576500:00011:00015",
  "USGS:05576900:00011:00001",
  "USGS:01010000:00011:00005",
  "USGS:01010000:00011:00030",
  "USGS:01010000:00011:00018",
  "USGS:01010000:00011:00026",
  "USGS:01010000:00011:00006",
  "USGS:01010000:00011:00008",
  "USGS:01010070:00011:00017",
  "USGS:01010070:00011:00018",
  "USGS:01010070:00011:00004",
  "USGS:01010070:00011:00002",
  "USGS:01010500:00011:00018",
  "USGS:01010500:00011:00025",
  "USGS:01010500:00011:00005",
  "USGS:01010500:00011:00002",
  "USGS:01011000:00011:00004",
  "USGS:05487980:00011:00007",
  "USGS:05488110:00011:00002",
  "USGS:05488110:00011:00001",
  "USGS:05488200:00011:00001",
  "USGS:05488200:00011:00003",
  "USGS:05488500:00011:00001",
  "USGS:05488500:00011:00003",
  "USGS:05489000:00011:00001",
  "USGS:05489000:00011:00003",
  "USGS:05489500:00011:00001",
  "USGS:05489500:00011:00003",
  "USGS:05490500:00011:00001",
  "USGS:05490500:00011:00003",
  "USGS:05494300:00011:00001",
  "USGS:05494300:00011:00002",
  "USGS:06483290:00011:00002",
  "USGS:06483290:00011:00001",
  "USGS:06483495:00011:00001",
  "USGS:06483500:00011:00001",
  "USGS:06483500:00011:00002",
  "USGS:06485500:00011:00001",
  "USGS:06485500:00011:00006",
  "USGS:06485500:00011:00022",
  "USGS:06599900:00011:00006",
  "USGS:06599900:00011:00001",
  "USGS:06599900:00011:00007",
  "USGS:06599950:00011:00004",
  "USGS:06600000:00011:00004",
  "USGS:06600030:00011:00001",
  "USGS:06600100:00011:00001",
  "USGS:06600100:00011:00002",
  "USGS:06600500:00011:00001",
  "USGS:06600500:00011:00002",
  "USGS:06602020:00011:00005",
  "USGS:06602020:00011:00001",
  "USGS:06602020:00011:00022",
  "USGS:06602400:00011:00001",
  "USGS:06602400:00011:00002",
  "USGS:06604000:00011:00017",
  "USGS:06604000:00011:00003",
  "USGS:06604200:00011:00015",
  "USGS:06604200:00011:00012",
  "USGS:06604440:00011:00012",
  "USGS:06604440:00011:00001",
  "USGS:06604440:00011:00002",
  "USGS:06604440:00011:00014",
  "USGS:06605000:00011:00001",
  "USGS:06605000:00011:00013",
  "USGS:06605750:00011:00001",
  "USGS:06605850:00011:00005",
  "USGS:06605850:00011:00002",
  "USGS:06606600:00011:00001",
  "USGS:06606600:00011:00002",
  "USGS:06607200:00011:00001",
  "USGS:06607200:00011:00002",
  "USGS:06607500:00011:00001",
  "USGS:06607500:00011:00002",
  "USGS:06608500:00011:00004",
  "USGS:06608500:00011:00001",
  "USGS:06608500:00011:00002",
  "USGS:06609500:00011:00001",
  "USGS:06609500:00011:00002",
  "USGS:06609560:00011:00003",
  "USGS:06610505:00011:00004",
  "USGS:06610505:00011:00002",
  "USGS:06610505:00011:00005",
  "USGS:06610505:00011:00006",
  "USGS:06610505:00011:00007",
  "USGS:06610505:00011:00008",
  "USGS:06805850:00011:00003",
  "USGS:06805850:00011:00001",
  "USGS:06805850:00011:00002",
  "USGS:06807410:00011:00001",
  "USGS:06807410:00011:00002",
  "USGS:06808500:00011:00001",
  "USGS:06808500:00011:00022",
  "USGS:06808820:00011:00003",
  "USGS:06808820:00011:00001",
  "USGS:06808820:00011:00002",
  "USGS:06809210:00011:00001",
  "USGS:06809210:00011:00002",
  "USGS:06809500:00011:00002",
  "USGS:06809500:00011:00026",
  "USGS:06809900:00011:00003",
  "USGS:06809900:00011:00001",
  "USGS:06809900:00011:00002",
  "USGS:06810000:00011:00001",
  "USGS:06810000:00011:00002",
  "USGS:06811800:00011:00001",
  "USGS:03252300:00011:00013",
  "USGS:02492100:00011:00001",
  "USGS:02492100:00011:00014",
  "USGS:02492111:00011:00013",
  "USGS:02492111:00011:00001",
  "USGS:02492511:00011:00001",
  "USGS:02492519:00011:00003",
  "USGS:02492519:00011:00001",
  "USGS:02492519:00011:00014",
  "USGS:02492600:00011:00004",
  "USGS:02492600:00011:00015",
  "USGS:06811875:00011:00001",
  "USGS:06817000:00011:00011",
  "USGS:06817000:00011:00012",
  "USGS:06817000:00011:00002",
  "USGS:06817000:00011:00019",
  "USGS:06817000:00011:00010",
  "USGS:06819185:00011:00001",
  "USGS:06819185:00011:00004",
  "USGS:06856600:00011:00001",
  "USGS:06856600:00011:00002",
  "USGS:06857050:00011:00013",
  "USGS:06857050:00011:00001",
  "USGS:06857100:00011:00004",
  "USGS:06857100:00011:00003",
  "USGS:06860000:00011:00004",
  "USGS:06860000:00011:00003",
  "USGS:06861000:00011:00004",
  "USGS:06861000:00011:00003",
  "USGS:06861500:00011:00004",
  "USGS:06861500:00011:00002",
  "USGS:06862700:00011:00004",
  "USGS:06862850:00011:00004",
  "USGS:06862850:00011:00003",
  "USGS:06863000:00011:00003",
  "USGS:06863000:00011:00002",
  "USGS:06863420:00011:00002",
  "USGS:06863420:00011:00001",
  "USGS:06863500:00011:00004",
  "USGS:06863500:00011:00003",
  "USGS:06864000:00011:00001",
  "USGS:06864000:00011:00002",
  "USGS:06864500:00011:00001",
  "USGS:06864500:00011:00002",
  "USGS:06865000:00011:00013",
  "USGS:06865000:00011:00001",
  "USGS:06865500:00011:00004",
  "USGS:06865500:00011:00003",
  "USGS:06866000:00011:00001",
  "USGS:06866000:00011:00003",
  "USGS:06866500:00011:00001",
  "USGS:06866500:00011:00002",
  "USGS:06866900:00011:00008",
  "USGS:06866900:00011:00007",
  "USGS:06867000:00011:00001",
  "USGS:06867000:00011:00002",
  "USGS:06898000:00011:00002",
  "USGS:06898000:00011:00018",
  "USGS:06903400:00011:00006",
  "USGS:06903400:00011:00002",
  "USGS:06903700:00011:00004",
  "USGS:06903700:00011:00002",
  "USGS:06903880:00011:00002",
  "USGS:06903900:00011:00002",
  "USGS:06903900:00011:00010",
  "USGS:06904010:00011:00005",
  "USGS:06904010:00011:00002",
  "USGS:404629095500501:00011:00001",
  "USCE:404753091054200:00011:00001",
  "USGS:410057095075101:00011:00001",
  "USGS:411843092105101:00011:00001",
  "USCE:412522091021200:00011:00001",
  "USGS:414315091252002:00011:00002",
  "USGS:415501096081201:00011:00001",
  "USGS:420117092505601:00011:00001",
  "USGS:421115091250501:00011:00001",
  "USCE:421539090252100:00011:00001",
  "USGS:430159093403201:00011:00001",
  "USGS:03288110:00011:00002",
  "USGS:03288110:00011:00001",
  "USGS:03288180:00011:00003",
  "USGS:03288180:00011:00002",
  "USGS:03288180:00011:00001",
  "USGS:03288190:00011:00002",
  "USGS:03288190:00011:00001",
  "USGS:03289000:00011:00005",
  "USGS:03289000:00011:00002",
  "USGS:03289000:00011:00004",
  "USGS:03289000:00011:00019",
  "USGS:03289000:00011:00022",
  "USGS:03289000:00011:00021",
  "USGS:402558087351501:00011:00001",
  "USCE:402715089362200:00011:00001",
  "USCE:402924090202500:00011:00001",
  "USCE:403725089143000:00011:00001",
  "USGS:404038089315201:00011:00002",
  "USGS:404038089315201:00011:00005",
  "USGS:404038089315201:00011:00003",
  "USGS:404038089315201:00011:00004",
  "USGS:404038089315201:00011:00001",
  "USGS:404038089315201:00011:00006",
  "USCE:404228090164800:00011:00001",
  "USCE:405240088381000:00011:00001",
  "USCE:405256091012600:00011:00001",
  "USCE:410005090511500:00011:00001",
  "USCE:410744090550900:00011:00001",
  "USCE:411113090580200:00011:00001",
  "USCE:411130091032900:00011:00001",
  "USCE:411230088555100:00011:00001",
  "USGS:411759088365101:00011:00005",
  "USGS:411759088365101:00011:00007",
  "USGS:411759088365101:00011:00004",
  "USGS:411759088365101:00011:00003",
  "USGS:411759088365101:00011:00001",
  "USGS:411759088365101:00011:00006",
  "USGS:411959088280101:00011:00015",
  "USGS:411959088280101:00011:00004",
  "USGS:411959088280101:00011:00003",
  "USGS:411959088280101:00011:00008",
  "USGS:411959088280101:00011:00009",
  "USGS:411959088280101:00011:00010",
  "USGS:411959088280101:00011:00011",
  "USGS:411959088280101:00011:00014",
  "USGS:411959088280101:00011:00012",
  "USGS:411959088280101:00011:00005",
  "USGS:411959088280101:00011:00013",
  "USGS:412033088264601:00011:00004",
  "USGS:412033088264601:00011:00006",
  "USGS:412033088264601:00011:00007",
  "USGS:412033088264601:00011:00008",
  "USGS:412033088264601:00011:00005",
  "USCE:412048088111100:00011:00001",
  "USGS:412104087573401:00011:00002",
  "USCE:412157089295400:00011:00001",
  "USGS:412320088154101:00011:00001",
  "USGS:412320088154101:00011:00004",
  "USGS:412354087370001:00011:00001",
  "USGS:412404088084801:00011:00002",
  "USGS:412429087504201:00011:00002",
  "USGS:412538087594301:00011:00002",
  "USGS:412657087372001:00011:00001",
  "USCE:412920090092700:00011:00001",
  "USGS:413102087510901:00011:00002",
  "USCE:413102090340000:00011:00001",
  "USGS:413113087342201:00011:00001",
  "USGS:413222087555101:00011:00002",
  "USCE:413322090110700:00011:00001",
  "USGS:413653087581901:00011:00002",
  "USGS:413718087440001:00011:00002",
  "USGS:413743089310101:00011:00001",
  "USGS:413743089310102:00011:00001",
  "USGS:414020088014601:00011:00006",
  "USGS:414020088014601:00011:00008",
  "USGS:414020088014601:00011:00004",
  "USGS:414020088014601:00011:00005",
  "USGS:414020088014601:00011:00003",
  "USGS:414020088014601:00011:00002",
  "USGS:414020088014601:00011:00007",
  "USGS:414205088193801:00011:00001",
  "USGS:414652088133800:00011:00004",
  "USCE:414658089445900:00011:00001",
  "USGS:414702088104801:00011:00002",
  "USGS:414903088101701:00011:00001",
  "USCE:414920087491500:00011:00001",
  "USGS:415037087581700:00011:00003",
  "USGS:03305000:00011:00001",
  "USGS:03305000:00011:00002",
  "USGS:03305990:00011:00002",
  "USGS:03305990:00011:00001",
  "USGS:03306000:00011:00003",
  "USGS:03306000:00011:00002",
  "USGS:03306500:00011:00001",
  "USGS:03306500:00011:00014",
  "USGS:03306500:00011:00004",
  "USGS:03307000:00011:00015",
  "USGS:03307000:00011:00004",
  "USGS:03307000:00011:00002",
  "USGS:07141000:00011:00002",
  "USGS:07141200:00011:00004",
  "USGS:07141200:00011:00003",
  "USGS:07141220:00011:00002",
  "USGS:07141220:00011:00001",
  "USGS:07141300:00011:00001",
  "USGS:07141300:00011:00002",
  "USGS:07141780:00011:00004",
  "USGS:07141780:00011:00003",
  "USGS:07141900:00011:00007",
  "USGS:07141900:00011:00006",
  "USGS:07142019:00011:00002",
  "USGS:07142019:00011:00001",
  "USGS:07142300:00011:00004",
  "USGS:07142300:00011:00003",
  "USGS:07142575:00011:00004",
  "USGS:07142575:00011:00003",
  "USGS:07142680:00011:00004",
  "USGS:07142680:00011:00003",
  "USGS:07143300:00011:00001",
  "USGS:07143300:00011:00002",
  "USGS:07143310:00011:00001",
  "USGS:07143330:00011:00001",
  "USGS:07143330:00011:00002",
  "USGS:07143375:00011:00005",
  "USGS:07143375:00011:00004",
  "USGS:07143665:00011:00004",
  "USGS:07143665:00011:00003",
  "USGS:07143672:00011:00016",
  "USGS:07143672:00011:00002",
  "USGS:07143672:00011:00001",
  "USGS:07143672:00011:00018",
  "USGS:07143672:00011:00019",
  "USGS:07143672:00011:00030",
  "USGS:07143672:00011:00033",
  "USGS:07143672:00011:00017",
  "USGS:07143672:00011:00020",
  "USGS:07143672:00011:00027",
  "USGS:07143672:00011:00029",
  "USGS:07144100:00011:00027",
  "USGS:07144100:00011:00054",
  "USGS:07144100:00011:00002",
  "USGS:07144100:00011:00001",
  "USGS:07144100:00011:00049",
  "USGS:07144100:00011:00029",
  "USGS:07144100:00011:00053",
  "USGS:07144100:00011:00030",
  "USGS:07144100:00011:00047",
  "USGS:07144100:00011:00056",
  "USGS:07144100:00011:00051",
  "USGS:07144100:00011:00057",
  "USGS:07144100:00011:00028",
  "USGS:07144100:00011:00055",
  "USGS:07144100:00011:00101",
  "USGS:07144100:00011:00052",
  "USGS:07144100:00011:00031",
  "USGS:07144100:00011:00044",
  "USGS:07144100:00011:00058",
  "USGS:07144100:00011:00064",
  "USGS:07144100:00011:00065",
  "USGS:07144100:00011:00046",
  "USGS:07144200:00011:00007",
  "USGS:07144200:00011:00006",
  "USGS:07144200:00011:00030",
  "USGS:07144201:00011:00002",
  "USGS:07144300:00011:00006",
  "USGS:07144300:00011:00005",
  "USGS:07144301:00011:00002",
  "USGS:07144301:00011:00001",
  "USGS:07144470:00011:00002",
  "USGS:07144480:00011:00001",
  "USGS:07144480:00011:00003",
  "USGS:07144480:00011:00002",
  "USGS:07144486:00011:00001",
  "USGS:07144486:00011:00002",
  "USGS:07144490:00011:00001",
  "USGS:07144490:00011:00002",
  "USGS:07144550:00011:00001",
  "USGS:07144550:00011:00002",
  "USGS:07144570:00011:00002",
  "USGS:07144570:00011:00001",
  "USGS:07144780:00011:00015",
  "USGS:07144780:00011:00004",
  "USGS:07144780:00011:00003",
  "USGS:07144780:00011:00016",
  "USGS:07144780:00011:00021",
  "USGS:07144780:00011:00030",
  "USGS:07144780:00011:00018",
  "USGS:07144780:00011:00023",
  "USGS:07144790:00011:00014",
  "USGS:07144790:00011:00029",
  "USGS:07144790:00011:00055",
  "USGS:07144790:00011:00056",
  "USGS:07144790:00011:00025",
  "USGS:07144790:00011:00017",
  "USGS:07144790:00011:00032",
  "USGS:07144790:00011:00057",
  "USGS:07144790:00011:00059",
  "USGS:07144790:00011:00016",
  "USGS:07144790:00011:00031",
  "USGS:07144790:00011:00021",
  "USGS:07144790:00011:00001",
  "USGS:07144790:00011:00024",
  "USGS:07144790:00011:00058",
  "USGS:07144790:00011:00064",
  "USGS:07144790:00011:00028",
  "USGS:07144795:00011:00004",
  "USGS:07144795:00011:00003",
  "USGS:07144910:00011:00004",
  "USGS:07144910:00011:00003",
  "USGS:07145200:00011:00001",
  "USGS:07145200:00011:00002",
  "USGS:07145500:00011:00001",
  "USGS:07145500:00011:00002",
  "USGS:07145600:00011:00011",
  "USGS:07145600:00011:00001",
  "USGS:07145700:00011:00004",
  "USGS:07145700:00011:00003",
  "USGS:07146500:00011:00001",
  "USGS:07146500:00011:00002",
  "USGS:07146800:00011:00002",
  "USGS:07146800:00011:00001",
  "USGS:07147070:00011:00001",
  "USGS:07147070:00011:00002",
  "USGS:07147190:00011:00001",
  "USGS:07147800:00011:00001",
  "USGS:07147800:00011:00002",
  "USGS:07147900:00011:00003",
  "USGS:07148111:00011:00002",
  "USGS:07148111:00011:00001",
  "USGS:07149000:00011:00012",
  "USGS:07149000:00011:00011",
  "USGS:07151500:00011:00007",
  "USGS:07151500:00011:00006",
  "USGS:07156900:00011:00005",
  "USGS:07156900:00011:00016",
  "USGS:07156900:00011:00015",
  "USGS:01021480:00011:00014",
  "USGS:01021480:00011:00015",
  "USGS:01021480:00011:00002",
  "USGS:01021480:00011:00001",
  "USGS:01022294:00011:00002",
  "USGS:01022294:00011:00001",
  "USGS:01022500:00011:00001",
  "USGS:01022500:00011:00023",
  "USGS:01022500:00011:00019",
  "USGS:01022500:00011:00021",
  "USGS:01022500:00011:00002",
  "USGS:01022500:00011:00006",
  "USGS:01022840:00011:00002",
  "USGS:01022840:00011:00001",
  "USGS:06876070:00011:00003",
  "USGS:06876440:00011:00001",
  "USGS:06876440:00011:00002",
  "USGS:06876700:00011:00004",
  "USGS:06876700:00011:00003",
  "USGS:06876900:00011:00001",
  "USGS:06876900:00011:00002",
  "USGS:06877600:00011:00001",
  "USGS:06877600:00011:00002",
  "USGS:06878000:00011:00006",
  "USGS:06878000:00011:00005",
  "USGS:06878600:00011:00003",
  "USGS:06878600:00011:00002",
  "USGS:06879100:00011:00001",
  "USGS:06879100:00011:00002",
  "USGS:06879100:00011:00016",
  "USGS:06879650:00011:00006",
  "USGS:06879650:00011:00005",
  "USGS:06879805:00011:00001",
  "USGS:06879810:00011:00002",
  "USGS:06879810:00011:00001",
  "USGS:06879815:00011:00001",
  "USGS:06879820:00011:00001",
  "USGS:06882510:00011:00001",
  "USGS:06882510:00011:00002",
  "USGS:06884025:00011:00006",
  "USGS:06884025:00011:00005",
  "USGS:06884200:00011:00004",
  "USGS:06884200:00011:00003",
  "USGS:06884400:00011:00001",
  "USGS:06884400:00011:00002",
  "USGS:06884700:00011:00001",
  "USGS:06885500:00011:00001",
  "USGS:06885500:00011:00002",
  "USGS:06886900:00011:00013",
  "USGS:06886900:00011:00001",
  "USGS:06887000:00011:00006",
  "USGS:06887000:00011:00005",
  "USGS:06887500:00011:00021",
  "USGS:06887500:00011:00039",
  "USGS:06887500:00011:00001",
  "USGS:06887500:00011:00002",
  "USGS:06887500:00011:00023",
  "USGS:06887500:00011:00040",
  "USGS:06887500:00011:00024",
  "USGS:06887500:00011:00043",
  "USGS:06887500:00011:00044",
  "USGS:06887500:00011:00022",
  "USGS:06887500:00011:00041",
  "USGS:06887500:00011:00045",
  "USGS:06887500:00011:00047",
  "USGS:06887500:00011:00029",
  "USGS:06887500:00011:00032",
  "USGS:06887500:00011:00042",
  "USGS:06887500:00011:00035",
  "USGS:06888000:00011:00006",
  "USGS:06888000:00011:00005",
  "USGS:06888350:00011:00014",
  "USGS:06888350:00011:00004",
  "USGS:06888350:00011:00003",
  "USGS:06888500:00011:00004",
  "USGS:06888500:00011:00003",
  "USGS:06888700:00011:00001",
  "USGS:06889000:00011:00001",
  "USGS:06889000:00011:00002",
  "USGS:06889200:00011:00004",
  "USGS:06889200:00011:00003",
  "USGS:06889500:00011:00004",
  "USGS:06889500:00011:00003",
  "USGS:06889585:00011:00001",
  "USGS:06889630:00011:00002",
  "USGS:06889630:00011:00001",
  "USGS:06890100:00011:00001",
  "USGS:06890100:00011:00002",
  "USGS:06890898:00011:00013",
  "USGS:06890898:00011:00001",
  "USGS:06890900:00011:00014",
  "USGS:06890900:00011:00017",
  "USGS:06890900:00011:00016",
  "USGS:06891000:00011:00001",
  "USGS:06891000:00011:00002",
  "USGS:01017290:00011:00002",
  "USGS:01017290:00011:00001",
  "USGS:01017550:00011:00002",
  "USGS:01017550:00011:00001",
  "USGS:01017960:00011:00002",
  "USGS:01017960:00011:00001",
  "USGS:01018000:00011:00001",
  "USGS:01018000:00011:00002",
  "USGS:01018009:00011:00002",
  "USGS:01018009:00011:00001",
  "USGS:01018035:00011:00012",
  "USGS:01495000:00011:00004",
  "USGS:07179300:00011:00001",
  "USGS:07179500:00011:00001",
  "USGS:07179500:00011:00002",
  "USGS:07179700:00011:00002",
  "USGS:07179700:00011:00001",
  "USGS:07179710:00011:00002",
  "USGS:07179730:00011:00001",
  "USGS:07179730:00011:00002",
  "USGS:07179750:00011:00002",
  "USGS:07179750:00011:00001",
  "USGS:07179795:00011:00001",
  "USGS:07179795:00011:00002",
  "USGS:07180200:00011:00002",
  "USGS:07180400:00011:00028",
  "USGS:07180400:00011:00002",
  "USGS:07180500:00011:00004",
  "USGS:07180500:00011:00003",
  "USGS:07182200:00011:00002",
  "USGS:07182200:00011:00001",
  "USGS:07182250:00011:00001",
  "USGS:07182250:00011:00002",
  "USGS:07182260:00011:00001",
  "USGS:07182260:00011:00002",
  "USGS:07182390:00011:00003",
  "USGS:07182390:00011:00002",
  "USGS:07182390:00011:00001",
  "USGS:07182390:00011:00004",
  "USGS:07182390:00011:00005",
  "USGS:07182510:00011:00016",
  "USGS:07182510:00011:00001",
  "USGS:07182510:00011:00002",
  "USGS:07182510:00011:00017",
  "USGS:07182510:00011:00018",
  "USGS:07183000:00011:00019",
  "USGS:07183000:00011:00001",
  "USGS:07183000:00011:00002",
  "USGS:07183000:00011:00020",
  "USGS:07183000:00011:00021",
  "USGS:07183300:00011:00001",
  "USGS:07183500:00011:00005",
  "USGS:07183500:00011:00001",
  "USGS:07183500:00011:00002",
  "USGS:07183500:00011:00007",
  "USGS:07183500:00011:00020",
  "USGS:07184000:00011:00004",
  "USGS:07184000:00011:00003",
  "USGS:07184500:00011:00001",
  "USGS:07184500:00011:00002",
  "USGS:07186055:00011:00002",
  "USGS:07186055:00011:00001",
  "USGS:07187600:00011:00001",
  "USGS:07187600:00011:00002",
  "USGS:370033100534202:00011:00001",
  "USGS:370033100534204:00011:00001",
  "USGS:370130101180902:00011:00001",
  "USGS:370130101180903:00011:00001",
  "USGS:374956097231601:00011:00001",
  "USGS:375259097252901:00011:00001",
  "USGS:375327097285401:00011:00003",
  "USGS:375327097285401:00011:00018",
  "USGS:375327097285401:00011:00007",
  "USGS:375327097285401:00011:00022",
  "USGS:375327097285401:00011:00002",
  "USGS:375327097285401:00011:00017",
  "USGS:375327097285401:00011:00005",
  "USGS:375327097285401:00011:00020",
  "USGS:375327097285401:00011:00006",
  "USGS:375327097285401:00011:00021",
  "USGS:375327097285401:00011:00004",
  "USGS:375327097285401:00011:00019",
  "USGS:375327097285401:00011:00023",
  "USGS:375327097285401:00011:00001",
  "USGS:375327097285402:00011:00003",
  "USGS:375327097285402:00011:00002",
  "USGS:375327097285402:00011:00005",
  "USGS:375327097285402:00011:00004",
  "USGS:375327097285402:00011:00001",
  "USGS:375332097284801:00011:00003",
  "USGS:375332097284801:00011:00018",
  "USGS:375332097284801:00011:00007",
  "USGS:375332097284801:00011:00022",
  "USGS:375332097284801:00011:00002",
  "USGS:375332097284801:00011:00017",
  "USGS:375332097284801:00011:00005",
  "USGS:375332097284801:00011:00020",
  "USGS:375332097284801:00011:00006",
  "USGS:375332097284801:00011:00021",
  "USGS:375332097284801:00011:00004",
  "USGS:375332097284801:00011:00019",
  "USGS:375332097284801:00011:00023",
  "USGS:375332097284801:00011:00001",
  "USGS:375332097284802:00011:00003",
  "USGS:375332097284802:00011:00002",
  "USGS:375332097284802:00011:00005",
  "USGS:375332097284802:00011:00004",
  "USGS:375332097284802:00011:00001",
  "USGS:375350097262800:00011:00012",
  "USGS:375350097262800:00011:00001",
  "USGS:375350097262800:00011:00011",
  "USGS:375350097262800:00011:00014",
  "USGS:375350097262800:00011:00015",
  "USGS:375350097262800:00011:00013",
  "USGS:375350097262800:00011:00017",
  "USGS:375350097262800:00011:00016",
  "USGS:375350097262800:00011:00018",
  "USGS:375642097385304:00011:00001",
  "USGS:375642097385305:00011:00001",
  "USGS:375814097324701:00011:00001",
  "USGS:375814097324702:00011:00001",
  "USGS:375936102023901:00011:00012",
  "USGS:375936102023901:00011:00011",
  "USGS:375936102023901:00011:00001",
  "USGS:01069700:00011:00001",
  "USGS:01069700:00011:00002",
  "USGS:06892350:00011:00001",
  "USGS:06892350:00011:00002",
  "USGS:06892350:00011:00020",
  "USGS:06892350:00011:00065",
  "USGS:06892350:00011:00021",
  "USGS:06892350:00011:00067",
  "USGS:06892350:00011:00068",
  "USGS:06892350:00011:00019",
  "USGS:06892350:00011:00066",
  "USGS:06892350:00011:00074",
  "USGS:06892350:00011:00071",
  "USGS:06892350:00011:00072",
  "USGS:06892350:00011:00025",
  "USGS:06892350:00011:00030",
  "USGS:06892350:00011:00069",
  "USGS:06892350:00011:00086",
  "USGS:06892360:00011:00002",
  "USGS:06892360:00011:00001",
  "USGS:06892493:00011:00001",
  "USGS:06892494:00011:00001",
  "USGS:06892495:00011:00004",
  "USGS:06892495:00011:00003",
  "USGS:06892513:00011:00027",
  "USGS:06892513:00011:00004",
  "USGS:06892513:00011:00003",
  "USGS:06892513:00011:00026",
  "USGS:06892513:00011:00029",
  "USGS:06892513:00011:00031",
  "USGS:06892513:00011:00028",
  "USGS:06892513:00011:00030",
  "USGS:06892950:00011:00001",
  "USGS:06893080:00011:00004",
  "USGS:06893080:00011:00003",
  "USGS:06893100:00011:00002",
  "USGS:06893100:00011:00001",
  "USGS:06893300:00011:00018",
  "USGS:06893300:00011:00001",
  "USGS:06893300:00011:00002",
  "USGS:06893300:00011:00017",
  "USGS:06893300:00011:00020",
  "USGS:06893300:00011:00019",
  "USGS:06893300:00011:00021",
  "USGS:06893350:00011:00013",
  "USGS:06893350:00011:00001",
  "USGS:06893350:00011:00002",
  "USGS:06893350:00011:00012",
  "USGS:06893350:00011:00015",
  "USGS:06893350:00011:00014",
  "USGS:06893350:00011:00016",
  "USGS:06893390:00011:00013",
  "USGS:06893390:00011:00054",
  "USGS:06893390:00011:00003",
  "USGS:06893390:00011:00002",
  "USGS:06893390:00011:00015",
  "USGS:06893390:00011:00053",
  "USGS:06893390:00011:00018",
  "USGS:06893390:00011:00056",
  "USGS:06893390:00011:00058",
  "USGS:06893390:00011:00014",
  "USGS:06893390:00011:00055",
  "USGS:06893390:00011:00016",
  "USGS:06893390:00011:00057",
  "USGS:06893390:00011:00052",
  "USGS:06893390:00011:00023",
  "USGS:06910800:00011:00001",
  "USGS:06910800:00011:00002",
  "USGS:06910997:00011:00013",
  "USGS:06910997:00011:00001",
  "USGS:06911000:00011:00001",
  "USGS:06911000:00011:00002",
  "USGS:06911490:00011:00006",
  "USGS:06911490:00011:00005",
  "USGS:06911900:00011:00004",
  "USGS:06911900:00011:00003",
  "USGS:06912490:00011:00013",
  "USGS:06912490:00011:00001",
  "USGS:06912500:00011:00004",
  "USGS:06912500:00011:00003",
  "USGS:06913000:00011:00004",
  "USGS:06913000:00011:00003",
  "USGS:06913500:00011:00001",
  "USGS:06913500:00011:00002",
  "USGS:06914100:00011:00002",
  "USGS:06914100:00011:00001",
  "USGS:06914500:00011:00001",
  "USGS:06914500:00011:00002",
  "USGS:06914950:00011:00002",
  "USGS:06914950:00011:00001",
  "USGS:06914990:00011:00002",
  "USGS:06914990:00011:00001",
  "USGS:06914995:00011:00013",
  "USGS:06914995:00011:00001",
  "USGS:06915000:00011:00001",
  "USGS:06915000:00011:00002",
  "USGS:06915800:00011:00001",
  "USGS:06915800:00011:00002",
  "USGS:06916600:00011:00001",
  "USGS:06916600:00011:00002",
  "USGS:06917000:00011:00004",
  "USGS:06917000:00011:00003",
  "USGS:06917240:00011:00002",
  "USGS:06917240:00011:00001",
  "USGS:06917500:00011:00001",
  "USGS:06917500:00011:00002",
  "USGS:07137000:00011:00001",
  "USGS:07137000:00011:00002",
  "USGS:07137000:00011:00006",
  "USGS:07137500:00011:00004",
  "USGS:07137500:00011:00001",
  "USGS:07137500:00011:00002",
  "USGS:07137500:00011:00006",
  "USGS:07138000:00011:00004",
  "USGS:07138000:00011:00003",
  "USGS:07138020:00011:00003",
  "USGS:07138020:00011:00002",
  "USGS:07138050:00011:00002",
  "USGS:07138050:00011:00001",
  "USGS:07138050:00011:00015",
  "USGS:07138063:00011:00002",
  "USGS:07138063:00011:00001",
  "USGS:07138063:00011:00015",
  "USGS:07138064:00011:00002",
  "USGS:07138064:00011:00001",
  "USGS:07138070:00011:00002",
  "USGS:07138070:00011:00001",
  "USGS:07138075:00011:00002",
  "USGS:07138075:00011:00001",
  "USGS:07138075:00011:00015",
  "USGS:07139000:00011:00004",
  "USGS:07139000:00011:00003",
  "USGS:07139500:00011:00005",
  "USGS:01581830:00011:00002",
  "USGS:01581830:00011:00001",
  "USGS:01581870:00011:00002",
  "USGS:01581870:00011:00001",
  "USGS:01581920:00011:00003",
  "USGS:01581920:00011:00002",
  "USGS:01581920:00011:00001",
  "USGS:01581960:00011:00002",
  "USGS:01581960:00011:00001",
  "USGS:01582000:00011:00001",
  "USGS:01582000:00011:00002",
  "USGS:01582500:00011:00001",
  "USGS:01582500:00011:00002",
  "USGS:01583100:00011:00001",
  "USGS:01583100:00011:00002",
  "USGS:01583500:00011:00001",
  "USGS:01583500:00011:00002",
  "USGS:01583570:00011:00001",
  "USGS:01583570:00011:00002",
  "USGS:01583580:00011:00002",
  "USGS:01027200:00011:00014",
  "USGS:01027200:00011:00015",
  "USGS:01027200:00011:00002",
  "USGS:01027200:00011:00001",
  "USGS:01029200:00011:00014",
  "USGS:01029200:00011:00015",
  "USGS:01029200:00011:00002",
  "USGS:01029200:00011:00001",
  "USGS:01029500:00011:00016",
  "USGS:01029500:00011:00017",
  "USGS:01029500:00011:00001",
  "USGS:01029500:00011:00002",
  "USGS:01030350:00011:00002",
  "USGS:01030350:00011:00001",
  "USGS:01030500:00011:00015",
  "USGS:01030500:00011:00017",
  "USGS:01030500:00011:00001",
  "USGS:01030500:00011:00003",
  "USGS:01031300:00011:00016",
  "USGS:01031300:00011:00018",
  "USGS:01031300:00011:00002",
  "USGS:01031300:00011:00001",
  "USGS:01031450:00011:00016",
  "USGS:01031450:00011:00018",
  "USGS:01031450:00011:00002",
  "USGS:01031450:00011:00001",
  "USGS:01031500:00011:00013",
  "USGS:01031500:00011:00027",
  "USGS:01031500:00011:00023",
  "USGS:01031500:00011:00024",
  "USGS:01031500:00011:00004",
  "USGS:01031500:00011:00002",
  "USGS:01031510:00011:00002",
  "USGS:01031510:00011:00001",
  "USGS:01034000:00011:00001",
  "USGS:01034000:00011:00002",
  "USGS:01034500:00011:00022",
  "USGS:01034500:00011:00023",
  "USGS:01034500:00011:00002",
  "USGS:01034500:00011:00006",
  "USGS:01036390:00011:00001",
  "USGS:01036390:00011:00039",
  "USGS:01036390:00011:00008",
  "USGS:01036390:00011:00003",
  "USGS:01036390:00011:00004",
  "USGS:01036390:00011:00029",
  "USGS:01036390:00011:00005",
  "USGS:01036390:00011:00031",
  "USGS:01037000:00011:00001",
  "USGS:01037000:00011:00002",
  "USGS:01037050:00011:00011",
  "USGS:01037380:00011:00016",
  "USGS:01037380:00011:00017",
  "USGS:01037380:00011:00014",
  "USGS:01037380:00011:00015",
  "USGS:01037380:00011:00002",
  "USGS:01037380:00011:00001",
  "USGS:01038000:00011:00001",
  "USGS:01038000:00011:00021",
  "USGS:01038000:00011:00018",
  "USGS:01038000:00011:00019",
  "USGS:01038000:00011:00002",
  "USGS:01038000:00011:00005",
  "USGS:01042500:00011:00020",
  "USGS:01042500:00011:00017",
  "USGS:01042500:00011:00001",
  "USGS:01042500:00011:00003",
  "USGS:01043500:00011:00001",
  "USGS:01043500:00011:00002",
  "USGS:01044550:00011:00017",
  "USGS:01044550:00011:00018",
  "USGS:01044550:00011:00002",
  "USGS:01044550:00011:00016",
  "USGS:01046000:00011:00001",
  "USGS:01046000:00011:00002",
  "USGS:01046500:00011:00023",
  "USGS:01046500:00011:00019",
  "USGS:01046500:00011:00002",
  "USGS:01046500:00011:00006",
  "USGS:01047000:00011:00022",
  "USGS:01047000:00011:00018",
  "USGS:01047000:00011:00004",
  "USGS:01047000:00011:00002",
  "USGS:01047150:00011:00002",
  "USGS:01047150:00011:00001",
  "USGS:01047200:00011:00002",
  "USGS:01047200:00011:00001",
  "USGS:01048000:00011:00019",
  "USGS:01048000:00011:00015",
  "USGS:01048000:00011:00002",
  "USGS:01048000:00011:00003",
  "USGS:01048220:00011:00002",
  "USGS:01048220:00011:00001",
  "USGS:01049265:00011:00004",
  "USGS:01049265:00011:00011",
  "USGS:01049320:00011:00001",
  "USGS:01049500:00011:00001",
  "USGS:01049500:00011:00003",
  "USGS:01049505:00011:00001",
  "USGS:01051715:00011:00001",
  "USGS:01054200:00011:00001",
  "USGS:01054200:00011:00023",
  "USGS:01054200:00011:00002",
  "USGS:01054200:00011:00004",
  "USGS:01054300:00011:00001",
  "USGS:01054300:00011:00002",
  "USGS:01054500:00011:00004",
  "USGS:01054500:00011:00002",
  "USGS:01055000:00011:00016",
  "USGS:01055000:00011:00017",
  "USGS:01055000:00011:00001",
  "USGS:01055000:00011:00003",
  "USGS:01055220:00011:00001",
  "USGS:01055500:00011:00001",
  "USGS:01055500:00011:00003",
  "USGS:01057000:00011:00020",
  "USGS:01057000:00011:00021",
  "USGS:01057000:00011:00003",
  "USGS:01057000:00011:00018",
  "USGS:01059000:00011:00001",
  "USGS:01059000:00011:00003",
  "USGS:01063310:00011:00002",
  "USGS:01063310:00011:00003",
  "USGS:01063995:00011:00002",
  "USGS:01064118:00011:00005",
  "USGS:01066000:00011:00024",
  "USGS:01066000:00011:00020",
  "USGS:01066000:00011:00002",
  "USGS:01066000:00011:00007",
  "USGS:01067950:00011:00002",
  "USGS:01067950:00011:00001",
  "USGS:01068910:00011:00002",
  "USGS:01068910:00011:00001",
  "USGS:01069500:00011:00001",
  "USGS:01069500:00011:00002",
  "USGS:01591700:00011:00001",
  "USGS:01591700:00011:00002",
  "USGS:01592500:00011:00001",
  "USGS:01592500:00011:00002",
  "USGS:01593370:00011:00002",
  "USGS:01593370:00011:00001",
  "USGS:01593450:00011:00002",
  "USGS:01593450:00011:00001",
  "USGS:01593500:00011:00001",
  "USGS:01593500:00011:00002",
  "USGS:01594000:00011:00001",
  "USGS:01594000:00011:00002",
  "USGS:01594440:00011:00002",
  "USGS:01594440:00011:00003",
  "USGS:01011000:00011:00019",
  "USGS:01011000:00011:00006",
  "USGS:01011000:00011:00002",
  "USGS:01013500:00011:00001",
  "USGS:01013500:00011:00021",
  "USGS:01014000:00011:00021",
  "USGS:01014000:00011:00022",
  "USGS:01014000:00011:00003",
  "USGS:01014000:00011:00019",
  "USGS:01015800:00011:00017",
  "USGS:01015800:00011:00020",
  "USGS:01015800:00011:00001",
  "USGS:01015800:00011:00023",
  "USGS:01017000:00011:00001",
  "USGS:01017000:00011:00005",
  "USGS:01017060:00011:00002",
  "USGS:01017060:00011:00001",
  "USGS:03213700:00011:00001",
  "USGS:03213700:00011:00003",
  "USGS:03215000:00011:00006",
  "USGS:03215410:00011:00012",
  "USGS:03215410:00011:00001",
  "USGS:03216000:00011:00001",
  "USGS:03216300:00011:00001",
  "USGS:03216350:00011:00004",
  "USGS:03216350:00011:00003",
  "USGS:03216350:00011:00002",
  "USGS:03216400:00011:00002",
  "USGS:03216500:00011:00003",
  "USGS:03216500:00011:00006",
  "USGS:03216500:00011:00002",
  "USGS:03216600:00011:00001",
  "USGS:03216600:00011:00018",
  "USGS:03217000:00011:00002",
  "USGS:03217000:00011:00003",
  "USGS:03238000:00011:00001",
  "USGS:03238140:00011:00003",
  "USGS:03238140:00011:00002",
  "USGS:03238140:00011:00001",
  "USGS:03238745:00011:00003",
  "USGS:03238745:00011:00002",
  "USGS:03238745:00011:00001",
  "USGS:03238772:00011:00003",
  "USGS:03238772:00011:00002",
  "USGS:03238772:00011:00001",
  "USGS:03248300:00011:00002",
  "USGS:03248300:00011:00001",
  "USGS:03249498:00011:00012",
  "USGS:03249498:00011:00002",
  "USGS:03249498:00011:00001",
  "USGS:03249500:00011:00002",
  "USGS:03249505:00011:00008",
  "USGS:03249505:00011:00007",
  "USGS:03250100:00011:00001",
  "USGS:03250100:00011:00002",
  "USGS:03250190:00011:00002",
  "USGS:03250190:00011:00001",
  "USGS:03250322:00011:00012",
  "USGS:03250322:00011:00002",
  "USGS:03250322:00011:00001",
  "USGS:03250500:00011:00001",
  "USGS:03250500:00011:00002",
  "USGS:03251200:00011:00013",
  "USGS:03251200:00011:00002",
  "USGS:03251200:00011:00001",
  "USGS:03251500:00011:00008",
  "USGS:03251500:00011:00002",
  "USGS:03251500:00011:00007",
  "USGS:375954097363801:00011:00003",
  "USGS:375954097363801:00011:00005",
  "USGS:375954097363801:00011:00001",
  "USGS:375954097363801:00011:00002",
  "USGS:375954097363801:00011:00016",
  "USGS:375954097363802:00011:00003",
  "USGS:375954097363802:00011:00005",
  "USGS:375954097363802:00011:00001",
  "USGS:375954097363802:00011:00002",
  "USGS:375954097363802:00011:00007",
  "USGS:380117102023801:00011:00012",
  "USGS:380117102023801:00011:00011",
  "USGS:380117102023801:00011:00001",
  "USGS:380643097353001:00011:00001",
  "USGS:381119098435301:00011:00001",
  "USGS:381421095451600:00011:00002",
  "USGS:381421095451600:00011:00001",
  "USGS:381421095451600:00011:00003",
  "USGS:384226099203801:00011:00001",
  "USGS:384242099165201:00011:00001",
  "USGS:03294570:00011:00016",
  "USGS:384253099180701:00011:00001",
  "USGS:384253099185201:00011:00001",
  "USGS:384259099195801:00011:00001",
  "USGS:390006095132301:00011:00001",
  "USGS:390601096433801:00011:00013",
  "USGS:390601096433801:00011:00003",
  "USGS:390644096430201:00011:00001",
  "USGS:390644096430202:00011:00001",
  "USGS:390823096455101:00011:00001",
  "USGS:390828096454706:00011:00002",
  "USGS:390828096454706:00011:00001",
  "USGS:04043238:00011:00011",
  "USGS:04043238:00011:00012",
  "USGS:04043238:00011:00010",
  "USGS:04043238:00011:00013",
  "USGS:04043244:00011:00003",
  "USGS:04043244:00011:00002",
  "USGS:04043244:00011:00001",
  "USGS:04043244:00011:00004",
  "USGS:04043275:00011:00012",
  "USGS:04043275:00011:00003",
  "USGS:04043275:00011:00001",
  "USGS:04043275:00011:00013",
  "USGS:04044724:00011:00002",
  "USGS:04044724:00011:00001",
  "USGS:04045500:00011:00001",
  "USGS:04045500:00011:00004",
  "USGS:04046000:00011:00002",
  "USGS:04046000:00011:00001",
  "USGS:01018035:00011:00020",
  "USGS:01018035:00011:00019",
  "USGS:01018035:00011:00002",
  "USGS:01018035:00011:00001",
  "USGS:01018035:00011:00021",
  "USGS:01018035:00011:00024",
  "USGS:01018035:00011:00023",
  "USGS:01018035:00011:00022",
  "USGS:01018500:00011:00001",
  "USGS:01018500:00011:00004",
  "USGS:01018900:00011:00002",
  "USGS:01018900:00011:00012",
  "USGS:01018900:00011:00001",
  "USGS:01019000:00011:00015",
  "USGS:01019000:00011:00017",
  "USGS:01019000:00011:00002",
  "USGS:01019000:00011:00001",
  "USGS:01019300:00011:00002",
  "USGS:01019300:00011:00012",
  "USGS:01019300:00011:00001",
  "USGS:01021000:00011:00004",
  "USGS:01021000:00011:00002",
  "USGS:01021470:00011:00002",
  "USGS:01021470:00011:00001",
  "USGS:0148471320:00011:00002",
  "USGS:0148471320:00011:00001",
  "USGS:01485000:00011:00001",
  "USGS:01485000:00011:00002",
  "USGS:01485500:00011:00001",
  "USGS:01485500:00011:00002",
  "USGS:01486000:00011:00001",
  "USGS:01486000:00011:00002",
  "USGS:01486500:00011:00001",
  "USGS:01486500:00011:00002",
  "USGS:01488110:00011:00001",
  "USGS:01490000:00011:00001",
  "USGS:01490000:00011:00002",
  "USGS:01491000:00011:00002",
  "USGS:01491000:00011:00003",
  "USGS:01491500:00011:00001",
  "USGS:01491500:00011:00002",
  "USGS:01492500:00011:00001",
  "USGS:01492500:00011:00002",
  "USGS:01493000:00011:00001",
  "USGS:01493000:00011:00002",
  "USGS:01493112:00011:00015",
  "USGS:01493112:00011:00002",
  "USGS:01493112:00011:00001",
  "USGS:01493112:00011:00016",
  "USGS:01493112:00011:00012",
  "USGS:01493112:00011:00010",
  "USGS:01493112:00011:00011",
  "USGS:01493112:00011:00014",
  "USGS:01493500:00011:00001",
  "USGS:01493500:00011:00002",
  "USGS:01494150:00011:00002",
  "USGS:01494150:00011:00001",
  "USGS:01495000:00011:00001",
  "USGS:01578310:00011:00002",
  "USGS:01578310:00011:00003",
  "USGS:01578475:00011:00002",
  "USGS:01578475:00011:00001",
  "USGS:01579550:00011:00001",
  "USGS:01579550:00011:00002",
  "USGS:01579550:00011:00005",
  "USGS:01579550:00011:00003",
  "USGS:01579550:00011:00006",
  "USGS:01579550:00011:00004",
  "USGS:01579550:00011:00008",
  "USGS:01580000:00011:00001",
  "USGS:01580000:00011:00002",
  "USGS:01580520:00011:00002",
  "USGS:01580520:00011:00001",
  "USGS:01580620:00011:00001",
  "USGS:01580620:00011:00003",
  "USGS:01580700:00011:00002",
  "USGS:01580700:00011:00001",
  "USGS:01581500:00011:00001",
  "USGS:01581500:00011:00002",
  "USGS:03437370:00011:00002",
  "USGS:03437370:00011:00001",
  "USGS:03437400:00011:00004",
  "USGS:03437400:00011:00001",
  "USGS:03437480:00011:00002",
  "USGS:03437480:00011:00003",
  "USGS:03437480:00011:00001",
  "USGS:03437495:00011:00002",
  "USGS:03437495:00011:00003",
  "USGS:03437495:00011:00001",
  "USGS:03437500:00011:00006",
  "USGS:03437500:00011:00002",
  "USGS:03437500:00011:00004",
  "USGS:03438000:00011:00003",
  "USGS:03438000:00011:00006",
  "USGS:03438000:00011:00002",
  "USGS:03610000:00011:00003",
  "USGS:03610000:00011:00001",
  "USGS:03610000:00011:00002",
  "USGS:03610200:00011:00001",
  "USGS:03610200:00011:00003",
  "USGS:03611000:00011:00002",
  "USGS:03611000:00011:00001",
  "USGS:07024000:00011:00002",
  "USGS:07024000:00011:00004",
  "USGS:365210088391301:00011:00003",
  "USGS:371954082350601:00011:00001",
  "USGS:372418082444201:00011:00001",
  "USGS:380249084295001:00011:00003",
  "USGS:381100082533601:00011:00001",
  "USGS:01646500:00011:00005",
  "USGS:01646500:00011:00006",
  "USGS:01646500:00011:00007",
  "USGS:01646500:00011:00022",
  "USGS:01646500:00011:00001",
  "USGS:01646500:00011:00002",
  "USGS:01646500:00011:00008",
  "USGS:01646500:00011:00023",
  "USGS:03289000:00011:00007",
  "USGS:03289193:00011:00005",
  "USGS:03289193:00011:00002",
  "USGS:03289193:00011:00001",
  "USGS:03289193:00011:00017",
  "USGS:03289193:00011:00019",
  "USGS:03289193:00011:00018",
  "USGS:03289200:00011:00003",
  "USGS:03289200:00011:00002",
  "USGS:03289200:00011:00001",
  "USGS:03289300:00011:00001",
  "USGS:03289300:00011:00002",
  "USGS:03289500:00011:00001",
  "USGS:03289500:00011:00002",
  "USGS:03289500:00011:00004",
  "USGS:03290080:00011:00011",
  "USGS:03290080:00011:00001",
  "USGS:03290080:00011:00013",
  "USGS:03290500:00011:00006",
  "USGS:03290500:00011:00002",
  "USGS:03291000:00011:00001",
  "USGS:03291000:00011:00002",
  "USGS:03291500:00011:00001",
  "USGS:03291500:00011:00002",
  "USGS:03292470:00011:00013",
  "USGS:03292470:00011:00002",
  "USGS:03292470:00011:00001",
  "USGS:03292470:00011:00017",
  "USGS:03292470:00011:00014",
  "USGS:03292470:00011:00016",
  "USGS:03292474:00011:00014",
  "USGS:03292474:00011:00002",
  "USGS:03292474:00011:00001",
  "USGS:03292474:00011:00018",
  "USGS:03292474:00011:00015",
  "USGS:03292474:00011:00017",
  "USGS:03292475:00011:00014",
  "USGS:03292475:00011:00002",
  "USGS:03292475:00011:00001",
  "USGS:03292475:00011:00017",
  "USGS:03292475:00011:00015",
  "USGS:03292475:00011:00018",
  "USGS:03292480:00011:00015",
  "USGS:03292480:00011:00002",
  "USGS:03292480:00011:00004",
  "USGS:03292480:00011:00018",
  "USGS:03292480:00011:00016",
  "USGS:03292480:00011:00019",
  "USGS:03292494:00011:00002",
  "USGS:03292494:00011:00001",
  "USGS:03292500:00011:00003",
  "USGS:03292500:00011:00001",
  "USGS:03292500:00011:00002",
  "USGS:03292500:00011:00004",
  "USGS:03292500:00011:00005",
  "USGS:03292500:00011:00006",
  "USGS:03292557:00011:00001",
  "USGS:03293000:00011:00003",
  "USGS:03293000:00011:00001",
  "USGS:03293000:00011:00002",
  "USGS:03293000:00011:00004",
  "USGS:03293000:00011:00005",
  "USGS:03293000:00011:00006",
  "USGS:03293500:00011:00003",
  "USGS:03293500:00011:00001",
  "USGS:03293500:00011:00008",
  "USGS:03293500:00011:00004",
  "USGS:03293500:00011:00005",
  "USGS:03293500:00011:00006",
  "USGS:03293510:00011:00002",
  "USGS:03293510:00011:00014",
  "USGS:03293510:00011:00016",
  "USGS:03293510:00011:00001",
  "USGS:03293510:00011:00018",
  "USGS:03293510:00011:00003",
  "USGS:03293510:00011:00017",
  "USGS:03293530:00011:00014",
  "USGS:03293530:00011:00002",
  "USGS:03293530:00011:00001",
  "USGS:03293530:00011:00019",
  "USGS:03293530:00011:00016",
  "USGS:03293530:00011:00018",
  "USGS:03294500:00011:00003",
  "USGS:03294500:00011:00002",
  "USGS:03294550:00011:00006",
  "USGS:03294550:00011:00005",
  "USGS:03294570:00011:00013",
  "USGS:03294570:00011:00002",
  "USGS:03294570:00011:00001",
  "USGS:03294570:00011:00014",
  "USGS:03294570:00011:00017",
  "USGS:03294600:00011:00001",
  "USGS:03295400:00011:00017",
  "USGS:03295400:00011:00002",
  "USGS:03295400:00011:00003",
  "USGS:03295597:00011:00014",
  "USGS:03295597:00011:00003",
  "USGS:03295597:00011:00004",
  "USGS:03295890:00011:00005",
  "USGS:03295890:00011:00001",
  "USGS:03295890:00011:00003",
  "USGS:03297800:00011:00013",
  "USGS:03297800:00011:00002",
  "USGS:03297800:00011:00001",
  "USGS:03297800:00011:00016",
  "USGS:03297800:00011:00014",
  "USGS:03297800:00011:00017",
  "USGS:03297900:00011:00015",
  "USGS:03297900:00011:00002",
  "USGS:03297900:00011:00003",
  "USGS:03297900:00011:00019",
  "USGS:03297900:00011:00016",
  "USGS:03297900:00011:00018",
  "USGS:03298000:00011:00015",
  "USGS:03298000:00011:00001",
  "USGS:03298000:00011:00002",
  "USGS:03298000:00011:00018",
  "USGS:03298000:00011:00016",
  "USGS:03298000:00011:00019",
  "USGS:03298135:00011:00018",
  "USGS:03298135:00011:00014",
  "USGS:03298135:00011:00016",
  "USGS:03298135:00011:00020",
  "USGS:03298135:00011:00021",
  "USGS:03298135:00011:00019",
  "USGS:03298150:00011:00007",
  "USGS:03298150:00011:00002",
  "USGS:03298150:00011:00005",
  "USGS:03298150:00011:00009",
  "USGS:03298150:00011:00010",
  "USGS:03298150:00011:00008",
  "USGS:03298200:00011:00015",
  "USGS:03298200:00011:00002",
  "USGS:03298200:00011:00001",
  "USGS:03298200:00011:00018",
  "USGS:03298200:00011:00016",
  "USGS:03298200:00011:00019",
  "USGS:03298250:00011:00015",
  "USGS:03298250:00011:00002",
  "USGS:03298250:00011:00001",
  "USGS:03298250:00011:00018",
  "USGS:03298250:00011:00016",
  "USGS:03298250:00011:00019",
  "USGS:03298300:00011:00016",
  "USGS:03298300:00011:00002",
  "USGS:03298300:00011:00005",
  "USGS:03298300:00011:00019",
  "USGS:03298300:00011:00017",
  "USGS:03298300:00011:00020",
  "USGS:03298470:00011:00001",
  "USGS:03298500:00011:00019",
  "USGS:03298500:00011:00005",
  "USGS:03298500:00011:00002",
  "USGS:03298550:00011:00011",
  "USGS:03298550:00011:00001",
  "USGS:03300400:00011:00018",
  "USGS:03300400:00011:00002",
  "USGS:03300400:00011:00003",
  "USGS:03301000:00011:00001",
  "USGS:03301000:00011:00002",
  "USGS:03301500:00011:00018",
  "USGS:03301500:00011:00005",
  "USGS:03301500:00011:00001",
  "USGS:03301630:00011:00001",
  "USGS:03301900:00011:00016",
  "USGS:03301900:00011:00002",
  "USGS:03301900:00011:00005",
  "USGS:03301900:00011:00019",
  "USGS:03301900:00011:00017",
  "USGS:03301900:00011:00020",
  "USGS:03301940:00011:00021",
  "USGS:03301940:00011:00001",
  "USGS:03301940:00011:00003",
  "USGS:03301940:00011:00024",
  "USGS:03301940:00011:00022",
  "USGS:03301940:00011:00025",
  "USGS:03302000:00011:00003",
  "USGS:03302000:00011:00001",
  "USGS:03302000:00011:00002",
  "USGS:03302000:00011:00004",
  "USGS:03302000:00011:00005",
  "USGS:03302000:00011:00006",
  "USGS:03302030:00011:00016",
  "USGS:03302030:00011:00002",
  "USGS:03302030:00011:00005",
  "USGS:03302030:00011:00019",
  "USGS:03302030:00011:00017",
  "USGS:03302030:00011:00020",
  "USGS:03302050:00011:00013",
  "USGS:03302050:00011:00002",
  "USGS:03302050:00011:00001",
  "USGS:03302050:00011:00017",
  "USGS:03302050:00011:00014",
  "USGS:03302050:00011:00016",
  "USGS:04108600:00011:00001",
  "USGS:04108600:00011:00002",
  "USGS:04108660:00011:00003",
  "USGS:04108660:00011:00002",
  "USGS:04108660:00011:00001",
  "USGS:04108660:00011:00007",
  "USGS:04108660:00011:00011",
  "USGS:04108660:00011:00008",
  "USGS:04108660:00011:00009",
  "USGS:04108800:00011:00001",
  "USGS:04108800:00011:00002",
  "USGS:04109000:00011:00001",
  "USGS:04109000:00011:00002",
  "USGS:04111000:00011:00001",
  "USGS:04111000:00011:00002",
  "USGS:04111379:00011:00001",
  "USGS:04111379:00011:00003",
  "USGS:04112000:00011:00001",
  "USGS:03252300:00011:00002",
  "USGS:03252300:00011:00001",
  "USGS:03252500:00011:00017",
  "USGS:03252500:00011:00002",
  "USGS:03253000:00011:00008",
  "USGS:03253000:00011:00004",
  "USGS:03253000:00011:00001",
  "USGS:03253000:00011:00002",
  "USGS:03253000:00011:00005",
  "USGS:03253500:00011:00004",
  "USGS:03253500:00011:00002",
  "USGS:03254480:00011:00003",
  "USGS:03254480:00011:00002",
  "USGS:03254480:00011:00001",
  "USGS:03254520:00011:00004",
  "USGS:03254520:00011:00003",
  "USGS:03254520:00011:00021",
  "USGS:03254520:00011:00002",
  "USGS:03254520:00011:00001",
  "USGS:03254520:00011:00008",
  "USGS:03254520:00011:00005",
  "USGS:03254520:00011:00007",
  "USGS:03254520:00011:00009",
  "USGS:03254520:00011:00026",
  "USGS:03254550:00011:00003",
  "USGS:03254550:00011:00002",
  "USGS:03254550:00011:00001",
  "USGS:03254693:00011:00003",
  "USGS:03254693:00011:00001",
  "USGS:03260015:00011:00003",
  "USGS:03260015:00011:00002",
  "USGS:03260015:00011:00001",
  "USGS:03260050:00011:00003",
  "USGS:03260050:00011:00002",
  "USGS:03260050:00011:00001",
  "USGS:03260100:00011:00003",
  "USGS:03260100:00011:00002",
  "USGS:03260100:00011:00001",
  "USGS:03262001:00011:00003",
  "USGS:03262001:00011:00002",
  "USGS:03262001:00011:00001",
  "USGS:03277075:00011:00013",
  "USGS:03277075:00011:00003",
  "USGS:03277075:00011:00002",
  "USGS:03277075:00011:00001",
  "USGS:03277075:00011:00017",
  "USGS:03277075:00011:00014",
  "USGS:03277075:00011:00016",
  "USGS:03277075:00011:00018",
  "USGS:03277130:00011:00004",
  "USGS:03277130:00011:00003",
  "USGS:03277130:00011:00002",
  "USGS:03277130:00011:00001",
  "USGS:03277130:00011:00008",
  "USGS:03277130:00011:00005",
  "USGS:03277130:00011:00007",
  "USGS:03277130:00011:00009",
  "USGS:03277200:00011:00008",
  "USGS:03277200:00011:00029",
  "USGS:03277200:00011:00034",
  "USGS:03277200:00011:00037",
  "USGS:03277200:00011:00002",
  "USGS:03277200:00011:00001",
  "USGS:03277200:00011:00012",
  "USGS:03277200:00011:00032",
  "USGS:03277200:00011:00035",
  "USGS:03277200:00011:00038",
  "USGS:03277200:00011:00030",
  "USGS:03277200:00011:00033",
  "USGS:03277200:00011:00036",
  "USGS:03277200:00011:00039",
  "USGS:03277200:00011:00040",
  "USGS:03277300:00011:00002",
  "USGS:03277300:00011:00013",
  "USGS:03277300:00011:00001",
  "USGS:03277446:00011:00003",
  "USGS:03277446:00011:00002",
  "USGS:03277446:00011:00001",
  "USGS:03277450:00011:00018",
  "USGS:03277450:00011:00002",
  "USGS:03277500:00011:00003",
  "USGS:03277500:00011:00002",
  "USGS:03280000:00011:00003",
  "USGS:03280000:00011:00006",
  "USGS:03280000:00011:00002",
  "USGS:03280600:00011:00016",
  "USGS:03280600:00011:00002",
  "USGS:03280700:00011:00003",
  "USGS:03280700:00011:00006",
  "USGS:03280700:00011:00002",
  "USGS:03280800:00011:00012",
  "USGS:03280800:00011:00002",
  "USGS:03280800:00011:00001",
  "USGS:03281000:00011:00020",
  "USGS:03281000:00011:00004",
  "USGS:03281000:00011:00002",
  "USGS:03281100:00011:00016",
  "USGS:03281100:00011:00001",
  "USGS:03281100:00011:00002",
  "USGS:03281500:00011:00020",
  "USGS:03281500:00011:00002",
  "USGS:03281500:00011:00006",
  "USGS:03282000:00011:00003",
  "USGS:03282000:00011:00005",
  "USGS:03282000:00011:00002",
  "USGS:03282040:00011:00002",
  "USGS:03282040:00011:00003",
  "USGS:03282060:00011:00011",
  "USGS:03282060:00011:00001",
  "USGS:03282120:00011:00002",
  "USGS:03282120:00011:00001",
  "USGS:03282290:00011:00002",
  "USGS:03282290:00011:00001",
  "USGS:03282500:00011:00001",
  "USGS:03282500:00011:00002",
  "USGS:03283500:00011:00005",
  "USGS:03283500:00011:00001",
  "USGS:03283500:00011:00003",
  "USGS:03284000:00011:00003",
  "USGS:03284000:00011:00006",
  "USGS:03284000:00011:00002",
  "USGS:03284230:00011:00002",
  "USGS:03284230:00011:00001",
  "USGS:03284500:00011:00002",
  "USGS:03284500:00011:00003",
  "USGS:03284525:00011:00003",
  "USGS:03284525:00011:00002",
  "USGS:03284525:00011:00001",
  "USGS:03284533:00011:00004",
  "USGS:03284533:00011:00002",
  "USGS:03284533:00011:00001",
  "USGS:03284552:00011:00004",
  "USGS:03284552:00011:00002",
  "USGS:03284552:00011:00001",
  "USGS:03284580:00011:00011",
  "USGS:03284580:00011:00001",
  "USGS:03285000:00011:00003",
  "USGS:03285000:00011:00006",
  "USGS:03285000:00011:00002",
  "USGS:03286000:00011:00001",
  "USGS:03286200:00011:00012",
  "USGS:03286200:00011:00002",
  "USGS:03286500:00011:00014",
  "USGS:03286500:00011:00002",
  "USGS:03286500:00011:00001",
  "USGS:03287000:00011:00005",
  "USGS:03287000:00011:00002",
  "USGS:03287000:00011:00006",
  "USGS:03287250:00011:00014",
  "USGS:03287250:00011:00001",
  "USGS:03287250:00011:00002",
  "USGS:03287500:00011:00001",
  "USGS:03287500:00011:00022",
  "USGS:03287500:00011:00002",
  "USGS:03287500:00011:00007",
  "USGS:03287590:00011:00003",
  "USGS:03287590:00011:00002",
  "USGS:03287590:00011:00001",
  "USGS:03287600:00011:00003",
  "USGS:03287600:00011:00002",
  "USGS:03287600:00011:00001",
  "USGS:03288100:00011:00002",
  "USGS:03288100:00011:00001",
  "USGS:04136500:00011:00004",
  "USGS:04136500:00011:00002",
  "USGS:04136500:00011:00001",
  "USGS:04136500:00011:00006",
  "USGS:04136900:00011:00004",
  "USGS:04136900:00011:00002",
  "USGS:04136900:00011:00003",
  "USGS:04136900:00011:00006",
  "USGS:04137005:00011:00003",
  "USGS:04137005:00011:00002",
  "USGS:04137005:00011:00001",
  "USGS:04137005:00011:00005",
  "USGS:04137020:00011:00001",
  "USGS:04137020:00011:00003",
  "USGS:04137025:00011:00001",
  "USGS:01094400:00011:00001",
  "USGS:01094400:00011:00003",
  "USGS:01094500:00011:00001",
  "USGS:01094500:00011:00002",
  "USGS:01095220:00011:00003",
  "USGS:01095220:00011:00008",
  "USGS:01095220:00011:00005",
  "USGS:01095220:00011:00002",
  "USGS:01095220:00011:00001",
  "USGS:01095220:00011:00004",
  "USGS:01095375:00011:00003",
  "USGS:01095375:00011:00006",
  "USGS:01095375:00011:00002",
  "USGS:01095375:00011:00001",
  "USGS:01095375:00011:00004",
  "USGS:01095434:00011:00007",
  "USGS:01095434:00011:00002",
  "USGS:01095434:00011:00001",
  "USGS:01095434:00011:00006",
  "USGS:01095503:00011:00012",
  "USGS:01095503:00011:00001",
  "USGS:01095503:00011:00002",
  "USGS:01095503:00011:00013",
  "USGS:01581649:00011:00002",
  "USGS:01581649:00011:00001",
  "USGS:01581700:00011:00001",
  "USGS:01581700:00011:00002",
  "USGS:01581752:00011:00004",
  "USGS:01581752:00011:00002",
  "USGS:01581752:00011:00001",
  "USGS:01581752:00011:00005",
  "USGS:01581752:00011:00006",
  "USGS:01581753:00011:00002",
  "USGS:01581753:00011:00001",
  "USGS:0158175320:00011:00002",
  "USGS:0158175320:00011:00001",
  "USGS:01581757:00011:00002",
  "USGS:01581757:00011:00001",
  "USGS:01581810:00011:00002",
  "USGS:01581810:00011:00001",
  "USGS:432310070393301:00011:00002",
  "USGS:434829070465101:00011:00003",
  "USGS:434955070261401:00011:00001",
  "USGS:435453070013601:00011:00001",
  "USGS:440213070203201:00011:00001",
  "USGS:440810069553601:00011:00001",
  "USGS:440823070291501:00011:00004",
  "USGS:440918069564001:00011:00001",
  "USGS:441801069455501:00011:00001",
  "USGS:441815069483401:00011:00002",
  "USGS:441815069483401:00011:00003",
  "USGS:441815069483401:00011:00001",
  "USGS:441815069483401:00011:00017",
  "USGS:442238068154101:00011:00001",
  "USGS:442450068175201:00011:00001",
  "USGS:443305070323701:00011:00002",
  "USGS:443305070323701:00011:00014",
  "USGS:443647070552303:00011:00001",
  "USGS:444227069561801:00011:00003",
  "USGS:444302070252401:00011:00001",
  "USGS:444950068220602:00011:00001",
  "USGS:445210069571901:00011:00003",
  "USGS:445227067520101:00011:00004",
  "USGS:445319068560101:00011:00004",
  "USGS:445810070463201:00011:00003",
  "USGS:445810070463201:00011:00004",
  "USGS:445810070463201:00011:00002",
  "USGS:450306069531101:00011:00002",
  "USGS:450306069531101:00011:00018",
  "USGS:450705069384801:00011:00001",
  "USGS:450705069384801:00011:00019",
  "USGS:450713067162801:00011:00001",
  "USGS:451031069185301:00011:00002",
  "USGS:451031069185301:00011:00017",
  "USGS:451105069270801:00011:00002",
  "USGS:451105069270801:00011:00004",
  "USGS:451317070115201:00011:00003",
  "USGS:451317070115201:00011:00004",
  "USGS:451317070115201:00011:00002",
  "USGS:451603069350101:00011:00002",
  "USGS:451603069350101:00011:00004",
  "USGS:452025069574701:00011:00003",
  "USGS:452156069371801:00011:00001",
  "USGS:452156069371801:00011:00016",
  "USGS:453405067254501:00011:00001",
  "USGS:453405067254501:00011:00005",
  "USGS:453629068531801:00011:00001",
  "USGS:463642069344601:00011:00004",
  "USGS:464200069425701:00011:00003",
  "USGS:470646069052501:00011:00002",
  "USGS:470646069052501:00011:00016",
  "USGS:471457068353001:00011:00004",
  "USGS:01096500:00011:00001",
  "USGS:01096500:00011:00003",
  "USGS:01097000:00011:00001",
  "USGS:01097000:00011:00005",
  "USGS:01097300:00011:00003",
  "USGS:01097300:00011:00007",
  "USGS:01098499:00011:00002",
  "USGS:01098499:00011:00001",
  "USGS:01098500:00011:00001",
  "USGS:01098500:00011:00002",
  "USGS:01098530:00011:00001",
  "USGS:01098530:00011:00003",
  "USGS:01099500:00011:00001",
  "USGS:01099500:00011:00015",
  "USGS:01100000:00011:00002",
  "USGS:01100000:00011:00008",
  "USGS:01100500:00011:00001",
  "USGS:01100568:00011:00003",
  "USGS:01100568:00011:00002",
  "USGS:01100568:00011:00001",
  "USGS:01100600:00011:00001",
  "USGS:01100600:00011:00003",
  "USGS:01100627:00011:00012",
  "USGS:04174500:00011:00006",
  "USGS:03308500:00011:00004",
  "USGS:03308500:00011:00005",
  "USGS:03308500:00011:00002",
  "USGS:03310000:00011:00001",
  "USGS:03310000:00011:00002",
  "USGS:03310300:00011:00001",
  "USGS:03310300:00011:00002",
  "USGS:03310400:00011:00001",
  "USGS:03310400:00011:00002",
  "USGS:03310900:00011:00003",
  "USGS:03310900:00011:00002",
  "USGS:03310900:00011:00001",
  "USGS:03311000:00011:00003",
  "USGS:03311000:00011:00001",
  "USGS:03311500:00011:00004",
  "USGS:03311500:00011:00003",
  "USGS:03311500:00011:00002",
  "USGS:03312900:00011:00001",
  "USGS:03313000:00011:00017",
  "USGS:03313000:00011:00003",
  "USGS:03313000:00011:00002",
  "USGS:03313700:00011:00001",
  "USGS:03313700:00011:00004",
  "USGS:03314000:00011:00003",
  "USGS:03314000:00011:00005",
  "USGS:03314000:00011:00002",
  "USGS:03314500:00011:00003",
  "USGS:03314500:00011:00006",
  "USGS:03314500:00011:00002",
  "USGS:03315500:00011:00004",
  "USGS:03316500:00011:00001",
  "USGS:03316500:00011:00004",
  "USGS:03316645:00011:00005",
  "USGS:03318005:00011:00003",
  "USGS:03318005:00011:00002",
  "USGS:03318005:00011:00001",
  "USGS:03318010:00011:00003",
  "USGS:03318010:00011:00001",
  "USGS:03318800:00011:00002",
  "USGS:03319000:00011:00002",
  "USGS:03319885:00011:00007",
  "USGS:03319885:00011:00005",
  "USGS:03320000:00011:00003",
  "USGS:03320000:00011:00006",
  "USGS:03320000:00011:00002",
  "USGS:03320500:00011:00001",
  "USGS:03320500:00011:00004",
  "USGS:03321350:00011:00001",
  "USGS:03321350:00011:00002",
  "USGS:03321500:00011:00001",
  "USGS:03321500:00011:00005",
  "USGS:03321500:00011:00007",
  "USGS:03321500:00011:00013",
  "USGS:03321500:00011:00004",
  "USGS:03321500:00011:00003",
  "USGS:03321500:00011:00008",
  "USGS:03321500:00011:00009",
  "USGS:03321500:00011:00010",
  "USGS:03321500:00011:00012",
  "USGS:03322190:00011:00002",
  "USGS:03322190:00011:00001",
  "USGS:03322420:00011:00003",
  "USGS:03322420:00011:00002",
  "USGS:03381700:00011:00004",
  "USGS:03381700:00011:00003",
  "USGS:03381700:00011:00002",
  "USGS:03381700:00011:00015",
  "USGS:03383000:00011:00002",
  "USGS:03383000:00011:00007",
  "USGS:03384100:00011:00013",
  "USGS:03384100:00011:00003",
  "USGS:03400500:00011:00003",
  "USGS:03400500:00011:00005",
  "USGS:03400500:00011:00002",
  "USGS:03400986:00011:00003",
  "USGS:03400986:00011:00002",
  "USGS:03400986:00011:00001",
  "USGS:03401000:00011:00003",
  "USGS:03401000:00011:00006",
  "USGS:03401000:00011:00002",
  "USGS:03401385:00011:00003",
  "USGS:03401385:00011:00001",
  "USGS:03401385:00011:00002",
  "USGS:03401385:00011:00006",
  "USGS:03401385:00011:00004",
  "USGS:03401385:00011:00005",
  "USGS:03401385:00011:00007",
  "USGS:03402900:00011:00003",
  "USGS:03402900:00011:00002",
  "USGS:03403500:00011:00003",
  "USGS:03403500:00011:00002",
  "USGS:03403910:00011:00001",
  "USGS:03403910:00011:00006",
  "USGS:03404000:00011:00003",
  "USGS:03404000:00011:00005",
  "USGS:03404000:00011:00002",
  "USGS:03404500:00011:00011",
  "USGS:03404500:00011:00002",
  "USGS:03404820:00011:00003",
  "USGS:03404820:00011:00002",
  "USGS:03404900:00011:00008",
  "USGS:03404900:00011:00002",
  "USGS:03406500:00011:00003",
  "USGS:03406500:00011:00006",
  "USGS:03406500:00011:00002",
  "USGS:03407500:00011:00001",
  "USGS:03407500:00011:00002",
  "USGS:03410500:00011:00003",
  "USGS:03410500:00011:00012",
  "USGS:03410500:00011:00002",
  "USGS:03413200:00011:00003",
  "USGS:03413200:00011:00001",
  "USGS:03413200:00011:00013",
  "USGS:03414100:00011:00003",
  "USGS:03414100:00011:00006",
  "USGS:03414100:00011:00001",
  "USGS:01102000:00011:00001",
  "USGS:01102000:00011:00003",
  "USGS:01102345:00011:00002",
  "USGS:01102345:00011:00001",
  "USGS:01102500:00011:00045",
  "USGS:01646500:00011:00015",
  "USGS:01646500:00011:00021",
  "USGS:01646500:00011:00016",
  "USGS:01646500:00011:00020",
  "USGS:01646500:00011:00014",
  "USGS:01646500:00011:00017",
  "USGS:01646500:00011:00010",
  "USGS:01647850:00011:00002",
  "USGS:01647850:00011:00001",
  "USGS:01649150:00011:00002",
  "USGS:01649150:00011:00001",
  "USGS:01649190:00011:00005",
  "USGS:01649190:00011:00002",
  "USGS:01649190:00011:00001",
  "USGS:01649190:00011:00004",
  "USGS:01649190:00011:00006",
  "USGS:01649190:00011:00003",
  "USGS:01649190:00011:00007",
  "USGS:01649500:00011:00003",
  "USGS:01649500:00011:00001",
  "USGS:01649500:00011:00002",
  "USGS:01649500:00011:00006",
  "USGS:01649500:00011:00007",
  "USGS:01649500:00011:00005",
  "USGS:01649500:00011:00008",
  "USGS:01650500:00011:00001",
  "USGS:01650500:00011:00002",
  "USGS:01650800:00011:00008",
  "USGS:01650800:00011:00002",
  "USGS:01650800:00011:00001",
  "USGS:01650800:00011:00011",
  "USGS:01650800:00011:00012",
  "USGS:01650800:00011:00010",
  "USGS:01650800:00011:00013",
  "USGS:01651000:00011:00002",
  "USGS:01651000:00011:00003",
  "USGS:01653600:00011:00001",
  "USGS:01653600:00011:00002",
  "USGS:01658000:00011:00002",
  "USGS:01658000:00011:00005",
  "USGS:01660920:00011:00001",
  "USGS:01660920:00011:00002",
  "USGS:01661050:00011:00001",
  "USGS:01661050:00011:00002",
  "USGS:01661500:00011:00001",
  "USGS:01661500:00011:00002",
  "USGS:03075500:00011:00005",
  "USGS:03075500:00011:00001",
  "USGS:03075500:00011:00002",
  "USGS:03075905:00011:00002",
  "USGS:03075905:00011:00001",
  "USGS:03076100:00011:00002",
  "USGS:03076100:00011:00001",
  "USGS:03076500:00011:00004",
  "USGS:03076500:00011:00002",
  "USGS:03076500:00011:00003",
  "USGS:03076600:00011:00001",
  "USGS:03076600:00011:00002",
  "USGS:03076700:00011:00002",
  "USGS:03076700:00011:00001",
  "USGS:03076800:00011:00002",
  "USGS:03076800:00011:00001",
  "USGS:03078000:00011:00004",
  "USGS:03078000:00011:00001",
  "USGS:03078000:00011:00002",
  "USGS:04001000:00011:00003",
  "USGS:04001000:00011:00001",
  "USGS:04001000:00011:00002",
  "USGS:04031000:00011:00001",
  "USGS:04031000:00011:00002",
  "USGS:04032000:00011:00001",
  "USGS:04032000:00011:00002",
  "USGS:04033000:00011:00001",
  "USGS:04033000:00011:00002",
  "USGS:04033500:00011:00001",
  "USGS:04033500:00011:00002",
  "USGS:04035995:00011:00013",
  "USGS:04035995:00011:00002",
  "USGS:04035995:00011:00001",
  "USGS:04036000:00011:00001",
  "USGS:04036000:00011:00002",
  "USGS:04037400:00011:00001",
  "USGS:04037500:00011:00001",
  "USGS:04037500:00011:00002",
  "USGS:04040000:00011:00003",
  "USGS:04040000:00011:00004",
  "USGS:04040000:00011:00001",
  "USGS:04040000:00011:00002",
  "USGS:04040000:00011:00007",
  "USGS:04040000:00011:00012",
  "USGS:04040000:00011:00009",
  "USGS:04040000:00011:00010",
  "USGS:04040260:00011:00002",
  "USGS:04040304:00011:00002",
  "USGS:04040500:00011:00001",
  "USGS:04040500:00011:00002",
  "USGS:04041500:00011:00003",
  "USGS:04041500:00011:00001",
  "USGS:04041500:00011:00002",
  "USGS:04043016:00011:00002",
  "USGS:04043021:00011:00002",
  "USGS:04043050:00011:00004",
  "USGS:04043050:00011:00001",
  "USGS:04043050:00011:00002",
  "USGS:04043097:00011:00004",
  "USGS:04043097:00011:00002",
  "USGS:04043097:00011:00005",
  "USGS:04043150:00011:00002",
  "USGS:04043150:00011:00003",
  "USGS:04043150:00011:00001",
  "USGS:04043150:00011:00004",
  "USGS:381956076275301:00011:00001",
  "USGS:382407076260301:00011:00001",
  "USGS:383239076354201:00011:00001",
  "USGS:384333076394701:00011:00001",
  "USGS:391328077185901:00011:00001",
  "USGS:391407077174001:00011:00001",
  "USGS:392931076410301:00011:00001",
  "USGS:393126076244301:00011:00001",
  "USGS:394008077005601:00011:00001",
  "USGS:394050079180901:00011:00001",
  "USGS:01110500:00011:00001",
  "USGS:01110500:00011:00002",
  "USGS:01111200:00011:00001",
  "USGS:01111200:00011:00008",
  "USGS:01111212:00011:00002",
  "USGS:01111212:00011:00001",
  "USGS:01111230:00011:00001",
  "USGS:01111230:00011:00010",
  "USGS:01111230:00011:00008",
  "USGS:01111230:00011:00006",
  "USGS:01111230:00011:00002",
  "USGS:01111230:00011:00012",
  "USGS:01111230:00011:00009",
  "USGS:01123360:00011:00001",
  "USGS:01123360:00011:00008",
  "USGS:01123600:00011:00001",
  "USGS:01123600:00011:00006",
  "USGS:01124350:00011:00001",
  "USGS:01124350:00011:00005",
  "USGS:01124500:00011:00001",
  "USGS:01124500:00011:00005",
  "USGS:01125000:00011:00001",
  "USGS:01125000:00011:00018",
  "USGS:01125000:00011:00005",
  "USGS:01162000:00011:00001",
  "USGS:01162000:00011:00002",
  "USGS:01162500:00011:00001",
  "USGS:01162500:00011:00003",
  "USGS:01583580:00011:00003",
  "USGS:01583600:00011:00001",
  "USGS:01583600:00011:00002",
  "USGS:01583800:00011:00002",
  "USGS:01583800:00011:00001",
  "USGS:0158397967:00011:00002",
  "USGS:0158397967:00011:00001",
  "USGS:01584050:00011:00001",
  "USGS:01584050:00011:00002",
  "USGS:01584500:00011:00001",
  "USGS:01584500:00011:00002",
  "USGS:01585090:00011:00002",
  "USGS:01585090:00011:00001",
  "USGS:01585100:00011:00001",
  "USGS:01585100:00011:00002",
  "USGS:01585104:00011:00002",
  "USGS:01585104:00011:00001",
  "USGS:01585200:00011:00001",
  "USGS:01585200:00011:00002",
  "USGS:01585219:00011:00002",
  "USGS:01585219:00011:00001",
  "USGS:01585225:00011:00002",
  "USGS:01585225:00011:00001",
  "USGS:01585230:00011:00002",
  "USGS:01585230:00011:00001",
  "USGS:01585500:00011:00001",
  "USGS:01585500:00011:00002",
  "USGS:01586000:00011:00001",
  "USGS:01586000:00011:00002",
  "USGS:01586210:00011:00001",
  "USGS:01586210:00011:00002",
  "USGS:01586610:00011:00001",
  "USGS:01586610:00011:00002",
  "USGS:01589000:00011:00001",
  "USGS:01589000:00011:00002",
  "USGS:01589000:00011:00003",
  "USGS:01589025:00011:00002",
  "USGS:01589025:00011:00001",
  "USGS:01589025:00011:00003",
  "USGS:01589035:00011:00002",
  "USGS:01589035:00011:00001",
  "USGS:01589035:00011:00003",
  "USGS:01589100:00011:00001",
  "USGS:01589100:00011:00002",
  "USGS:01589180:00011:00002",
  "USGS:01589180:00011:00001",
  "USGS:01589197:00011:00002",
  "USGS:01589197:00011:00001",
  "USGS:01589238:00011:00002",
  "USGS:01589238:00011:00001",
  "USGS:01589290:00011:00002",
  "USGS:01589290:00011:00001",
  "USGS:01589300:00011:00002",
  "USGS:01589300:00011:00003",
  "USGS:01589305:00011:00002",
  "USGS:01589305:00011:00001",
  "USGS:01589312:00011:00002",
  "USGS:01589312:00011:00001",
  "USGS:01589315:00011:00001",
  "USGS:01589316:00011:00002",
  "USGS:01589316:00011:00001",
  "USGS:01589317:00011:00002",
  "USGS:01589317:00011:00001",
  "USGS:01589320:00011:00002",
  "USGS:01589320:00011:00001",
  "USGS:01589330:00011:00001",
  "USGS:01589330:00011:00002",
  "USGS:01589352:00011:00002",
  "USGS:01589352:00011:00001",
  "USGS:01589440:00011:00001",
  "USGS:01589440:00011:00002",
  "USGS:01589464:00011:00002",
  "USGS:01589464:00011:00001",
  "USGS:01589500:00011:00001",
  "USGS:01589500:00011:00002",
  "USGS:01589795:00011:00002",
  "USGS:01589795:00011:00001",
  "USGS:01591000:00011:00001",
  "USGS:01591000:00011:00002",
  "USGS:01591400:00011:00001",
  "USGS:01591400:00011:00002",
  "USGS:01591610:00011:00004",
  "USGS:01591610:00011:00001",
  "USGS:01591610:00011:00002",
  "USGS:02430085:00011:00004",
  "USGS:02430085:00011:00003",
  "USGS:02430680:00011:00004",
  "USGS:02430680:00011:00003",
  "USGS:02430880:00011:00004",
  "USGS:02430880:00011:00003",
  "USGS:01100627:00011:00013",
  "USGS:01100627:00011:00001",
  "USGS:01100627:00011:00002",
  "USGS:01100693:00011:00001",
  "USGS:01101000:00011:00001",
  "USGS:01101000:00011:00003",
  "USGS:01101500:00011:00001",
  "USGS:01101500:00011:00003",
  "USGS:04010500:00011:00019",
  "USGS:04010500:00011:00016",
  "USGS:04010500:00011:00015",
  "USGS:04010500:00011:00018",
  "USGS:04168580:00011:00002",
  "USGS:04168580:00011:00001",
  "USGS:04170000:00011:00001",
  "USGS:04170000:00011:00002",
  "USGS:04170500:00011:00001",
  "USGS:04170500:00011:00002",
  "USGS:04172000:00011:00001",
  "USGS:04172000:00011:00002",
  "USGS:04173500:00011:00001",
  "USGS:04173500:00011:00002",
  "USGS:04174490:00011:00004",
  "USGS:04174490:00011:00007",
  "USGS:04174490:00011:00002",
  "USGS:04174500:00011:00004",
  "USGS:04174500:00011:00001",
  "USGS:04174500:00011:00002",
  "USGS:04174500:00011:00007",
  "USGS:04174500:00011:00005",
  "USGS:04174500:00011:00018",
  "USGS:04174518:00011:00002",
  "USGS:04174518:00011:00001",
  "USGS:04175600:00011:00001",
  "USGS:04175600:00011:00002",
  "USGS:04176000:00011:00001",
  "USGS:04176000:00011:00002",
  "USGS:04176400:00011:00002",
  "USGS:04176500:00011:00006",
  "USGS:04176500:00011:00001",
  "USGS:04176500:00011:00004",
  "USGS:04176500:00011:00002",
  "USGS:04176500:00011:00008",
  "USGS:04176500:00011:00007",
  "USGS:04176500:00011:00010",
  "USGS:415318085243401:00011:00001",
  "USGS:415602084593701:00011:00001",
  "USGS:421332085401901:00011:00001",
  "USGS:421332085401902:00011:00001",
  "USGS:421435085353701:00011:00001",
  "USGS:421435085353702:00011:00001",
  "USGS:421448085383601:00011:00001",
  "USGS:421457085325801:00011:00001",
  "USGS:421614085270801:00011:00001",
  "USGS:421614085354001:00011:00001",
  "USGS:421641085350601:00011:00001",
  "USGS:421716085373702:00011:00001",
  "USGS:421918085283801:00011:00001",
  "USGS:422239083032401:00011:00005",
  "USGS:422239083032401:00011:00003",
  "USGS:422239083032401:00011:00004",
  "USGS:422239083032401:00011:00001",
  "USGS:422239083032401:00011:00006",
  "USGS:422239083032401:00011:00009",
  "USGS:422239083032401:00011:00007",
  "USGS:422517083131601:00011:00006",
  "USGS:422517083131601:00011:00003",
  "USGS:422517083131601:00011:00004",
  "USGS:422517083131601:00011:00001",
  "USGS:422517083131601:00011:00005",
  "USGS:422517083131601:00011:00010",
  "USGS:422517083131601:00011:00007",
  "USGS:422517083131601:00011:00008",
  "USGS:434103083130301:00011:00001",
  "USGS:442400084472801:00011:00001",
  "USGS:442409084274001:00011:00001",
  "USGS:442805084411001:00011:00001",
  "USGS:445512084415301:00011:00001",
  "USGS:450415085153501:00011:00001",
  "USGS:454427084424002:00011:00001",
  "USGS:05061000:00011:00007",
  "USGS:05061000:00011:00008",
  "USGS:05061000:00011:00010",
  "USGS:05061500:00011:00002",
  "USGS:05061500:00011:00007",
  "USGS:05061500:00011:00009",
  "USGS:05061500:00011:00019",
  "USGS:01594526:00011:00001",
  "USGS:01594526:00011:00002",
  "USGS:01594950:00011:00005",
  "USGS:01594950:00011:00004",
  "USGS:01594963:00011:00002",
  "USGS:01594963:00011:00001",
  "USGS:01595000:00011:00001",
  "USGS:01595000:00011:00002",
  "USGS:01595500:00011:00002",
  "USGS:01595500:00011:00003",
  "USGS:01595790:00011:00001",
  "USGS:01596050:00011:00002",
  "USGS:01596050:00011:00001",
  "USGS:01596500:00011:00006",
  "USGS:01596500:00011:00001",
  "USGS:01596500:00011:00002",
  "USGS:01597000:00011:00002",
  "USGS:01597000:00011:00003",
  "USGS:01597490:00011:00001",
  "USGS:01597500:00011:00005",
  "USGS:01597500:00011:00001",
  "USGS:01597500:00011:00002",
  "USGS:01598650:00011:00001",
  "USGS:01599000:00011:00002",
  "USGS:01599000:00011:00003",
  "USGS:01601100:00011:00002",
  "USGS:01601100:00011:00001",
  "USGS:01601500:00011:00001",
  "USGS:01601500:00011:00002",
  "USGS:01603000:00011:00002",
  "USGS:01603000:00011:00003",
  "USGS:01609000:00011:00001",
  "USGS:01609000:00011:00002",
  "USGS:01610000:00011:00002",
  "USGS:01610000:00011:00003",
  "USGS:01610155:00011:00001",
  "USGS:01610155:00011:00002",
  "USGS:01613000:00011:00002",
  "USGS:01613000:00011:00003",
  "USGS:01613095:00011:00002",
  "USGS:01613095:00011:00001",
  "USGS:01613525:00011:00002",
  "USGS:01613525:00011:00001",
  "USGS:01614500:00011:00002",
  "USGS:01614500:00011:00003",
  "USGS:01617800:00011:00001",
  "USGS:01617800:00011:00002",
  "USGS:01619000:00011:00001",
  "USGS:01619000:00011:00002",
  "USGS:01619500:00011:00002",
  "USGS:01619500:00011:00003",
  "USGS:01637500:00011:00002",
  "USGS:01637500:00011:00003",
  "USGS:01638500:00011:00002",
  "USGS:01638500:00011:00003",
  "USGS:01639000:00011:00001",
  "USGS:01639000:00011:00002",
  "USGS:01639500:00011:00001",
  "USGS:01639500:00011:00002",
  "USGS:01640975:00011:00001",
  "USGS:01642190:00011:00002",
  "USGS:01642190:00011:00001",
  "USGS:01643000:00011:00002",
  "USGS:01643000:00011:00003",
  "USGS:01643395:00011:00002",
  "USGS:01643395:00011:00001",
  "USGS:01643500:00011:00002",
  "USGS:01643500:00011:00003",
  "USGS:01644148:00011:00001",
  "USGS:01644371:00011:00002",
  "USGS:01644371:00011:00001",
  "USGS:01644372:00011:00002",
  "USGS:01644372:00011:00001",
  "USGS:01644375:00011:00002",
  "USGS:01644375:00011:00001",
  "USGS:01644380:00011:00002",
  "USGS:01644380:00011:00001",
  "USGS:01644388:00011:00002",
  "USGS:01644388:00011:00001",
  "USGS:01644390:00011:00002",
  "USGS:01644390:00011:00001",
  "USGS:01645000:00011:00001",
  "USGS:01645000:00011:00002",
  "USGS:05205900:00011:00001",
  "USGS:05207600:00011:00002",
  "USGS:05207600:00011:00001",
  "USGS:05210000:00011:00001",
  "USGS:05211000:00011:00012",
  "USGS:05211000:00011:00011",
  "USGS:05212700:00011:00001",
  "USGS:01102500:00011:00040",
  "USGS:01102500:00011:00026",
  "USGS:01102500:00011:00005",
  "USGS:01103025:00011:00003",
  "USGS:01103025:00011:00004",
  "USGS:01103025:00011:00001",
  "USGS:01103280:00011:00002",
  "USGS:01103280:00011:00003",
  "USGS:01103455:00011:00002",
  "USGS:01103500:00011:00005",
  "USGS:01103500:00011:00002",
  "USGS:01104000:00011:00001",
  "USGS:01104000:00011:00004",
  "USGS:01104200:00011:00001",
  "USGS:01104200:00011:00004",
  "USGS:01104370:00011:00004",
  "USGS:01104370:00011:00002",
  "USGS:01104370:00011:00001",
  "USGS:01104370:00011:00005",
  "USGS:01104405:00011:00003",
  "USGS:01104405:00011:00002",
  "USGS:01104405:00011:00001",
  "USGS:01104405:00011:00004",
  "USGS:01104415:00011:00003",
  "USGS:01104415:00011:00002",
  "USGS:01104415:00011:00001",
  "USGS:01104415:00011:00004",
  "USGS:01104415:00011:00019",
  "USGS:01104420:00011:00018",
  "USGS:01104420:00011:00001",
  "USGS:01104420:00011:00017",
  "USGS:01104430:00011:00003",
  "USGS:01104430:00011:00013",
  "USGS:01104430:00011:00014",
  "USGS:01104430:00011:00002",
  "USGS:01104430:00011:00011",
  "USGS:01104430:00011:00001",
  "USGS:01104430:00011:00004",
  "USGS:01104430:00011:00012",
  "USGS:01104430:00011:00030",
  "USGS:01104453:00011:00003",
  "USGS:01104453:00011:00002",
  "USGS:01104453:00011:00001",
  "USGS:01104453:00011:00004",
  "USGS:01104455:00011:00003",
  "USGS:01104455:00011:00002",
  "USGS:01104455:00011:00001",
  "USGS:01104455:00011:00004",
  "USGS:01104455:00011:00015",
  "USGS:01104455:00011:00023",
  "USGS:01104460:00011:00003",
  "USGS:01104460:00011:00002",
  "USGS:01104460:00011:00001",
  "USGS:01104460:00011:00004",
  "USGS:01104460:00011:00031",
  "USGS:01104475:00011:00003",
  "USGS:01104475:00011:00002",
  "USGS:01104475:00011:00001",
  "USGS:01104475:00011:00004",
  "USGS:01104475:00011:00019",
  "USGS:01104480:00011:00003",
  "USGS:01104480:00011:00010",
  "USGS:01104480:00011:00038",
  "USGS:01104480:00011:00039",
  "USGS:01104480:00011:00011",
  "USGS:01104480:00011:00002",
  "USGS:01104480:00011:00005",
  "USGS:01104480:00011:00001",
  "USGS:01104480:00011:00004",
  "USGS:01104480:00011:00013",
  "USGS:01104500:00011:00001",
  "USGS:01104500:00011:00003",
  "USGS:01104501:00011:00001",
  "USGS:01104501:00011:00002",
  "USGS:01104683:00011:00004",
  "USGS:01104683:00011:00001",
  "USGS:01104705:00011:00001",
  "USGS:01104715:00011:00001",
  "USGS:01104715:00011:00003",
  "USGS:01105000:00011:00001",
  "USGS:01105000:00011:00011",
  "USGS:01105500:00011:00001",
  "USGS:01105500:00011:00003",
  "USGS:01105554:00011:00002",
  "USGS:01105554:00011:00003",
  "USGS:011055566:00011:00003",
  "USGS:011055566:00011:00006",
  "USGS:01105583:00011:00002",
  "USGS:01105583:00011:00001",
  "USGS:01105584:00011:00002",
  "USGS:01105584:00011:00001",
  "USGS:01105585:00011:00004",
  "USGS:01105585:00011:00002",
  "USGS:01105600:00011:00001",
  "USGS:01105600:00011:00003",
  "USGS:01105606:00011:00004",
  "USGS:01105606:00011:00001",
  "USGS:01105607:00011:00003",
  "USGS:01105608:00011:00002",
  "USGS:01105608:00011:00001",
  "USGS:01105638:00011:00002",
  "USGS:01105730:00011:00002",
  "USGS:01105730:00011:00004",
  "USGS:01105870:00011:00002",
  "USGS:01105870:00011:00007",
  "USGS:01105876:00011:00002",
  "USGS:01105876:00011:00004",
  "USGS:01105880:00011:00001",
  "USGS:01105880:00011:00002",
  "USGS:011058837:00011:00002",
  "USGS:011058837:00011:00001",
  "USGS:01105933:00011:00002",
  "USGS:01105933:00011:00003",
  "USGS:01108000:00011:00001",
  "USGS:01108000:00011:00003",
  "USGS:01108410:00011:00002",
  "USGS:01108410:00011:00001",
  "USGS:01109000:00011:00001",
  "USGS:01109000:00011:00006",
  "USGS:01109060:00011:00001",
  "USGS:01109060:00011:00002",
  "USGS:01109070:00011:00001",
  "USGS:01109070:00011:00002",
  "USGS:01109730:00011:00001",
  "USGS:01109730:00011:00002",
  "USGS:01110000:00011:00001",
  "USGS:01110000:00011:00005",
  "USGS:07381343:00011:00006",
  "USGS:07381343:00011:00007",
  "USGS:07381343:00011:00005",
  "USGS:07381343:00011:00001",
  "USGS:07381343:00011:00003",
  "USGS:05338500:00011:00006",
  "USGS:05338500:00011:00005",
  "USGS:05341550:00011:00002",
  "USGS:05341550:00011:00014",
  "USGS:05341550:00011:00020",
  "USGS:05341550:00011:00013",
  "USGS:05341550:00011:00001",
  "USGS:05345000:00011:00012",
  "USGS:05345000:00011:00011",
  "USGS:05346050:00011:00001",
  "USGS:05346050:00011:00014",
  "USGS:05353800:00011:00009",
  "USGS:05353800:00011:00020",
  "USGS:05354500:00011:00001",
  "USGS:05355024:00011:00003",
  "USGS:05355024:00011:00002",
  "USGS:05355024:00011:00001",
  "USGS:02431000:00011:00005",
  "USGS:02431000:00011:00004",
  "USGS:02431000:00011:00003",
  "USGS:02432500:00011:00004",
  "USGS:02432500:00011:00003",
  "USGS:02433500:00011:00001",
  "USGS:02433500:00011:00020",
  "USGS:04015438:00011:00003",
  "USGS:04015438:00011:00002",
  "USGS:04015438:00011:00001",
  "USGS:04021520:00011:00002",
  "USGS:04021520:00011:00001",
  "USGS:04024000:00011:00001",
  "USGS:04024000:00011:00014",
  "USGS:04024000:00011:00006",
  "USGS:04024000:00011:00005",
  "USGS:04024000:00011:00004",
  "USGS:04024000:00011:00022",
  "USGS:04024000:00011:00023",
  "USGS:04024000:00011:00021",
  "USGS:04024000:00011:00024",
  "USGS:05030500:00011:00005",
  "USGS:05030500:00011:00015",
  "USGS:05046000:00011:00004",
  "USGS:05046000:00011:00003",
  "USGS:05046475:00011:00001",
  "USGS:05046475:00011:00002",
  "USGS:05049000:00011:00004",
  "USGS:05051300:00011:00002",
  "USGS:05051300:00011:00014",
  "USGS:413801070322703:00011:00001",
  "USGS:414100070011101:00011:00002",
  "USGS:414100070011101:00011:00001",
  "USGS:414124070265901:00011:00002",
  "USGS:414124070265901:00011:00001",
  "USGS:414124070311401:00011:00002",
  "USGS:414129070361401:00011:00002",
  "USGS:414129070361401:00011:00001",
  "USGS:414139070311501:00011:00002",
  "USGS:414159070310501:00011:00001",
  "USGS:414219070313601:00011:00002",
  "USGS:414630070014901:00011:00001",
  "USGS:414714071175901:00011:00002",
  "USGS:414714071175901:00011:00001",
  "USGS:415228070554601:00011:00001",
  "USGS:415353069585401:00011:00001",
  "USGS:415453070434901:00011:00002",
  "USGS:415453070434901:00011:00001",
  "USGS:420206070045901:00011:00002",
  "USGS:420206070045901:00011:00001",
  "USGS:420259072581701:00011:00003",
  "USGS:420259072581701:00011:00001",
  "USGS:420321070433502:00011:00001",
  "USGS:420351073193602:00011:00001",
  "USGS:420545071174001:00011:00001",
  "USGS:421852071220501:00011:00001",
  "USGS:422103072241102:00011:00004",
  "USGS:422103072241102:00011:00001",
  "USGS:422302071083801:00011:00002",
  "USGS:422302071083801:00011:00003",
  "USGS:422302071083801:00011:00005",
  "USGS:422302071083801:00011:00001",
  "USGS:422302071083801:00011:00004",
  "USGS:422302071083801:00011:00007",
  "USGS:422302071083801:00011:00006",
  "USGS:422328072035300:00011:00001",
  "USGS:422336072142100:00011:00002",
  "USGS:422341071464901:00011:00001",
  "USGS:422518071162501:00011:00002",
  "USGS:422518071162501:00011:00004",
  "USGS:422518071162501:00011:00005",
  "USGS:422518071162501:00011:00006",
  "USGS:422518071162501:00011:00008",
  "USGS:422518071162501:00011:00009",
  "USGS:422518071162501:00011:00012",
  "USGS:422518071162501:00011:00010",
  "USGS:422745073112001:00011:00001",
  "USGS:422812071244401:00011:00001",
  "USGS:422906072124301:00011:00001",
  "USGS:423115071032001:00011:00001",
  "USGS:423211071004400:00011:00002",
  "USGS:423401071093801:00011:00001",
  "USGS:423505070491702:00011:00002",
  "USGS:423505070491702:00011:00001",
  "USGS:423701071344800:00011:00002",
  "USGS:423815073100400:00011:00006",
  "USGS:423815073100400:00011:00008",
  "USGS:423815073100400:00011:00005",
  "USGS:423815073100400:00011:00004",
  "USGS:423815073100400:00011:00002",
  "USGS:423815073100400:00011:00007",
  "USGS:424520070562401:00011:00001",
  "USGS:424841071004101:00011:00001",
  "USGS:07344425:00011:00001",
  "USGS:07344425:00011:00013",
  "USGS:07344450:00011:00003",
  "USGS:07344460:00011:00001",
  "USGS:07344460:00011:00012",
  "USGS:07344480:00011:00001",
  "USGS:07346310:00011:00001",
  "USGS:07346450:00011:00001",
  "USGS:07346450:00011:00012",
  "USGS:07348000:00011:00007",
  "USGS:07348000:00011:00019",
  "USGS:07348098:00011:00001",
  "USGS:07348098:00011:00013",
  "USGS:07348500:00011:00005",
  "USGS:07348500:00011:00016",
  "USGS:07348550:00011:00001",
  "USGS:07348555:00011:00001",
  "USGS:07348700:00011:00006",
  "USGS:07348700:00011:00002",
  "USGS:07348700:00011:00005",
  "USGS:07349000:00011:00004",
  "USGS:07349250:00011:00001",
  "USGS:07349250:00011:00015",
  "USGS:07349298:00011:00001",
  "USGS:04056500:00011:00012",
  "USGS:04056500:00011:00001",
  "USGS:04056500:00011:00002",
  "USGS:04057510:00011:00001",
  "USGS:04057510:00011:00002",
  "USGS:04057800:00011:00004",
  "USGS:04057800:00011:00001",
  "USGS:04057800:00011:00003",
  "USGS:04057811:00011:00001",
  "USGS:04057812:00011:00002",
  "USGS:04057813:00011:00001",
  "USGS:04057813:00011:00003",
  "USGS:04057814:00011:00001",
  "USGS:04057814:00011:00003",
  "USGS:04058100:00011:00001",
  "USGS:04058100:00011:00002",
  "USGS:04058190:00011:00001",
  "USGS:04058200:00011:00001",
  "USGS:04058200:00011:00003",
  "USGS:04058940:00011:00001",
  "USGS:04059000:00011:00003",
  "USGS:04059000:00011:00005",
  "USGS:04059000:00011:00001",
  "USGS:04059000:00011:00004",
  "USGS:04059500:00011:00006",
  "USGS:04059500:00011:00001",
  "USGS:04059500:00011:00004",
  "USGS:04059500:00011:00003",
  "USGS:04059500:00011:00009",
  "USGS:04059500:00011:00007",
  "USGS:04059500:00011:00008",
  "USGS:04060500:00011:00001",
  "USGS:04060500:00011:00002",
  "USGS:04060993:00011:00002",
  "USGS:04060993:00011:00001",
  "USGS:04062000:00011:00001",
  "USGS:04062000:00011:00003",
  "USGS:04062500:00011:00001",
  "USGS:04062500:00011:00002",
  "USGS:04063500:00011:00002",
  "USGS:04063500:00011:00004",
  "USGS:04063500:00011:00001",
  "USGS:04063500:00011:00003",
  "USGS:04065650:00011:00002",
  "USGS:04065650:00011:00001",
  "USGS:04065722:00011:00002",
  "USGS:04065722:00011:00001",
  "USGS:04066003:00011:00005",
  "USGS:04066003:00011:00001",
  "USGS:04066003:00011:00002",
  "USGS:04066030:00011:00003",
  "USGS:04066030:00011:00008",
  "USGS:04066030:00011:00002",
  "USGS:04066030:00011:00004",
  "USGS:04066800:00011:00003",
  "USGS:04066800:00011:00002",
  "USGS:04066800:00011:00001",
  "USGS:04096015:00011:00002",
  "USGS:04096015:00011:00001",
  "USGS:04096405:00011:00002",
  "USGS:04096405:00011:00001",
  "USGS:04096515:00011:00001",
  "USGS:04096515:00011:00002",
  "USGS:04097188:00011:00001",
  "USGS:04097500:00011:00001",
  "USGS:04097500:00011:00002",
  "USGS:040975299:00011:00001",
  "USGS:040975299:00011:00002",
  "USGS:04097540:00011:00004",
  "USGS:04097540:00011:00001",
  "USGS:04097540:00011:00002",
  "USGS:04098980:00011:00001",
  "USGS:04098980:00011:00002",
  "USGS:04099000:00011:00001",
  "USGS:04099000:00011:00002",
  "USGS:04101500:00011:00003",
  "USGS:04101500:00011:00001",
  "USGS:04101500:00011:00004",
  "USGS:04101500:00011:00002",
  "USGS:04101500:00011:00006",
  "USGS:04101500:00011:00005",
  "USGS:04101500:00011:00009",
  "USGS:04101535:00011:00001",
  "USGS:04101535:00011:00002",
  "USGS:04101800:00011:00001",
  "USGS:04101800:00011:00002",
  "USGS:04102500:00011:00001",
  "USGS:04102500:00011:00002",
  "USGS:04102700:00011:00001",
  "USGS:04102700:00011:00002",
  "USGS:04103500:00011:00001",
  "USGS:04103500:00011:00002",
  "USGS:04104945:00011:00002",
  "USGS:04104945:00011:00001",
  "USGS:04105000:00011:00001",
  "USGS:04105000:00011:00002",
  "USGS:04105500:00011:00001",
  "USGS:04105500:00011:00002",
  "USGS:04105700:00011:00001",
  "USGS:04105700:00011:00002",
  "USGS:04106000:00011:00001",
  "USGS:04106000:00011:00002",
  "USGS:04106400:00011:00001",
  "USGS:04106400:00011:00002",
  "USGS:07369649:00011:00001",
  "USGS:07369700:00011:00002",
  "USGS:07369700:00011:00003",
  "USGS:07370000:00011:00005",
  "USGS:07371500:00011:00006",
  "USGS:07372050:00011:00002",
  "USGS:07372050:00011:00001",
  "USGS:07372190:00011:00001",
  "USGS:07372200:00011:00005",
  "USGS:07372200:00011:00013",
  "USGS:07373000:00011:00002",
  "USGS:07373000:00011:00004",
  "USGS:07374000:00011:00014",
  "USGS:07374000:00011:00022",
  "USGS:07374000:00011:00002",
  "USGS:05062000:00011:00008",
  "USGS:05062000:00011:00010",
  "USGS:05062500:00011:00002",
  "USGS:05062500:00011:00003",
  "USGS:05062500:00011:00022",
  "USGS:05063398:00011:00002",
  "USGS:05063398:00011:00001",
  "USGS:05063398:00011:00013",
  "USGS:05064000:00011:00006",
  "USGS:05064000:00011:00005",
  "USGS:05067500:00011:00004",
  "USGS:05067500:00011:00003",
  "USGS:05069000:00011:00001",
  "USGS:05069000:00011:00003",
  "USGS:05073500:00011:00001",
  "USGS:05073650:00011:00001",
  "USGS:05074000:00011:00003",
  "USGS:05074500:00011:00003",
  "USGS:05074500:00011:00004",
  "USGS:05075000:00011:00003",
  "USGS:05076000:00011:00004",
  "USGS:05076000:00011:00015",
  "USGS:05078000:00011:00006",
  "USGS:05078000:00011:00001",
  "USGS:05078230:00011:00001",
  "USGS:05078230:00011:00005",
  "USGS:05078470:00011:00004",
  "USGS:05078470:00011:00001",
  "USGS:05078500:00011:00001",
  "USGS:05078500:00011:00002",
  "USGS:05078500:00011:00004",
  "USGS:05078500:00011:00006",
  "USGS:05078520:00011:00004",
  "USGS:05078520:00011:00001",
  "USGS:05078720:00011:00002",
  "USGS:05078720:00011:00001",
  "USGS:05078770:00011:00004",
  "USGS:05078770:00011:00001",
  "USGS:05079000:00011:00006",
  "USGS:05079000:00011:00005",
  "USGS:05079200:00011:00004",
  "USGS:05079200:00011:00001",
  "USGS:05079250:00011:00004",
  "USGS:05079250:00011:00001",
  "USGS:05080000:00011:00002",
  "USGS:05080000:00011:00001",
  "USGS:05080000:00011:00013",
  "USGS:05083500:00011:00004",
  "USGS:05085450:00011:00002",
  "USGS:05085450:00011:00001",
  "USGS:05087500:00011:00002",
  "USGS:05087500:00011:00003",
  "USGS:05094000:00011:00005",
  "USGS:05094000:00011:00002",
  "USGS:05094000:00011:00004",
  "USGS:05104500:00011:00007",
  "USGS:05104500:00011:00001",
  "USGS:05104500:00011:00016",
  "USGS:05106000:00011:00001",
  "USGS:05106000:00011:00002",
  "USGS:05106000:00011:00013",
  "USGS:05107500:00011:00012",
  "USGS:05107500:00011:00004",
  "USGS:05107500:00011:00013",
  "USGS:05112000:00011:00006",
  "USGS:05112000:00011:00005",
  "USGS:05124480:00011:00001",
  "USGS:05124480:00011:00015",
  "USGS:05124480:00011:00008",
  "USGS:05124480:00011:00007",
  "USGS:05124982:00011:00002",
  "USGS:05124982:00011:00001",
  "USGS:05125000:00011:00013",
  "USGS:05125000:00011:00001",
  "USGS:05125000:00011:00002",
  "USGS:05125039:00011:00002",
  "USGS:05125039:00011:00001",
  "USGS:05126210:00011:00001",
  "USGS:05126210:00011:00002",
  "USGS:05127500:00011:00004",
  "USGS:05127500:00011:00003",
  "USGS:05129115:00011:00004",
  "USGS:05129115:00011:00003",
  "USGS:05129290:00011:00004",
  "USGS:05129290:00011:00003",
  "USGS:05129515:00011:00018",
  "USGS:05129515:00011:00014",
  "USGS:05129515:00011:00002",
  "USGS:05129515:00011:00019",
  "USGS:05129515:00011:00001",
  "USGS:05131500:00011:00021",
  "USGS:05131500:00011:00018",
  "USGS:05131500:00011:00008",
  "USGS:05131500:00011:00007",
  "USGS:05132000:00011:00006",
  "USGS:05132000:00011:00005",
  "USGS:05132000:00011:00002",
  "USGS:05132000:00011:00004",
  "USGS:05133500:00011:00001",
  "USGS:05133500:00011:00019",
  "USGS:05133500:00011:00006",
  "USGS:05133500:00011:00005",
  "USGS:05134200:00011:00003",
  "USGS:05134200:00011:00001",
  "USGS:05134200:00011:00002",
  "USGS:05134200:00011:00004",
  "USGS:05137500:00011:00003",
  "USGS:05137500:00011:00008",
  "USGS:05137500:00011:00002",
  "USGS:05137500:00011:00001",
  "USGS:05137500:00011:00004",
  "USGS:05140520:00011:00016",
  "USGS:05140520:00011:00004",
  "USGS:05140520:00011:00015",
  "USGS:05140521:00011:00003",
  "USGS:05200510:00011:00001",
  "USGS:05200510:00011:00004",
  "USGS:05200510:00011:00003",
  "USGS:07378500:00011:00006",
  "USGS:04137025:00011:00003",
  "USGS:04137030:00011:00001",
  "USGS:04137030:00011:00003",
  "USGS:04137500:00011:00003",
  "USGS:04137500:00011:00001",
  "USGS:04137500:00011:00004",
  "USGS:04137500:00011:00002",
  "USGS:04137500:00011:00007",
  "USGS:04137500:00011:00008",
  "USGS:04137500:00011:00009",
  "USGS:04142000:00011:00015",
  "USGS:04142000:00011:00002",
  "USGS:04142000:00011:00006",
  "USGS:04142000:00011:00001",
  "USGS:04142000:00011:00017",
  "USGS:04142000:00011:00018",
  "USGS:04142000:00011:00019",
  "USGS:04144500:00011:00001",
  "USGS:04144500:00011:00003",
  "USGS:04146000:00011:00001",
  "USGS:04146000:00011:00002",
  "USGS:04146063:00011:00001",
  "USGS:04146063:00011:00002",
  "USGS:04147500:00011:00001",
  "USGS:04147500:00011:00002",
  "USGS:04148140:00011:00001",
  "USGS:04148140:00011:00002",
  "USGS:0414826544:00011:00001",
  "USGS:0414826544:00011:00002",
  "USGS:0414826545:00011:00003",
  "USGS:0414826545:00011:00001",
  "USGS:0414826545:00011:00002",
  "USGS:0414826545:00011:00009",
  "USGS:0414826545:00011:00010",
  "USGS:041482663:00011:00006",
  "USGS:041482663:00011:00003",
  "USGS:041482663:00011:00001",
  "USGS:041482663:00011:00002",
  "USGS:041482663:00011:00008",
  "USGS:041482663:00011:00011",
  "USGS:041482663:00011:00009",
  "USGS:041482663:00011:00010",
  "USGS:04148300:00011:00002",
  "USGS:04148440:00011:00002",
  "USGS:04148500:00011:00001",
  "USGS:04148500:00011:00002",
  "USGS:04150800:00011:00002",
  "USGS:04151500:00011:00001",
  "USGS:04151500:00011:00002",
  "USGS:04152238:00011:00001",
  "USGS:04152238:00011:00002",
  "USGS:04152500:00011:00003",
  "USGS:04154000:00011:00001",
  "USGS:04154000:00011:00002",
  "USGS:04155500:00011:00002",
  "USGS:04155500:00011:00012",
  "USGS:04156000:00011:00001",
  "USGS:04156000:00011:00002",
  "USGS:04157005:00011:00001",
  "USGS:04157005:00011:00011",
  "USGS:04157005:00011:00009",
  "USGS:04157005:00011:00010",
  "USGS:04157005:00011:00003",
  "USGS:04157005:00011:00002",
  "USGS:04157005:00011:00006",
  "USGS:04157005:00011:00005",
  "USGS:04157060:00011:00005",
  "USGS:04157060:00011:00002",
  "USGS:04159010:00011:00002",
  "USGS:04159130:00011:00003",
  "USGS:04159130:00011:00004",
  "USGS:04159130:00011:00013",
  "USGS:04159492:00011:00002",
  "USGS:04159492:00011:00001",
  "USGS:04159900:00011:00001",
  "USGS:04159900:00011:00002",
  "USGS:04160600:00011:00001",
  "USGS:04160600:00011:00002",
  "USGS:04161000:00011:00001",
  "USGS:04161000:00011:00002",
  "USGS:04161540:00011:00001",
  "USGS:04161540:00011:00002",
  "USGS:04161820:00011:00001",
  "USGS:04161820:00011:00002",
  "USGS:04163400:00011:00001",
  "USGS:04163400:00011:00002",
  "USGS:04164000:00011:00001",
  "USGS:04164000:00011:00002",
  "USGS:04164100:00011:00001",
  "USGS:04164100:00011:00002",
  "USGS:04164300:00011:00002",
  "USGS:04164500:00011:00001",
  "USGS:04164500:00011:00002",
  "USGS:04164800:00011:00001",
  "USGS:04164800:00011:00002",
  "USGS:04165500:00011:00012",
  "USGS:04165500:00011:00011",
  "USGS:04165500:00011:00002",
  "USGS:04165500:00011:00001",
  "USGS:04165500:00011:00013",
  "USGS:04165500:00011:00016",
  "USGS:04165500:00011:00014",
  "USGS:04165500:00011:00015",
  "USGS:04165710:00011:00004",
  "USGS:04165710:00011:00001",
  "USGS:04165710:00011:00020",
  "USGS:04166000:00011:00001",
  "USGS:04166000:00011:00002",
  "USGS:04166100:00011:00001",
  "USGS:04166100:00011:00002",
  "USGS:04166300:00011:00001",
  "USGS:04166300:00011:00002",
  "USGS:04166500:00011:00003",
  "USGS:04166500:00011:00001",
  "USGS:04166500:00011:00002",
  "USGS:04166500:00011:00010",
  "USGS:04166500:00011:00006",
  "USGS:04166500:00011:00009",
  "USGS:04166500:00011:00011",
  "USGS:04167000:00011:00001",
  "USGS:04167000:00011:00002",
  "USGS:04168000:00011:00001",
  "USGS:04168000:00011:00002",
  "USGS:073814675:00011:00003",
  "USGS:073814675:00011:00002",
  "USGS:073814675:00011:00013",
  "USGS:073814675:00011:00001",
  "USGS:073814675:00011:00015",
  "USGS:073814675:00011:00017",
  "USGS:07381482:00011:00018",
  "USGS:07381482:00011:00003",
  "USGS:07381482:00011:00019",
  "USGS:07381482:00011:00001",
  "USGS:07381482:00011:00013",
  "USGS:07381490:00011:00020",
  "USGS:07381490:00011:00018",
  "USGS:07381495:00011:00003",
  "USGS:07381515:00011:00001",
  "USGS:073815450:00011:00001",
  "USGS:073815450:00011:00012",
  "USGS:07381567:00011:00013",
  "USGS:07381567:00011:00012",
  "USGS:07381567:00011:00001",
  "USGS:07381590:00011:00014",
  "USGS:07381590:00011:00024",
  "USGS:07381590:00011:00013",
  "USGS:073815925:00011:00001",
  "USGS:073815945:00011:00001",
  "USGS:073815963:00011:00002",
  "USGS:073815963:00011:00001",
  "USGS:04112000:00011:00002",
  "USGS:04112500:00011:00001",
  "USGS:04112500:00011:00002",
  "USGS:04112850:00011:00001",
  "USGS:04112850:00011:00002",
  "USGS:04113000:00011:00001",
  "USGS:04113000:00011:00002",
  "USGS:04114000:00011:00001",
  "USGS:04114000:00011:00004",
  "USGS:04114498:00011:00002",
  "USGS:04114498:00011:00001",
  "USGS:04115000:00011:00001",
  "USGS:04115000:00011:00002",
  "USGS:04115265:00011:00002",
  "USGS:04115265:00011:00001",
  "USGS:04116000:00011:00001",
  "USGS:04116000:00011:00002",
  "USGS:04116500:00011:00002",
  "USGS:04117000:00011:00001",
  "USGS:04117000:00011:00002",
  "USGS:04117500:00011:00001",
  "USGS:04117500:00011:00002",
  "USGS:04118000:00011:00002",
  "USGS:04118105:00011:00001",
  "USGS:04118500:00011:00001",
  "USGS:04118500:00011:00002",
  "USGS:04119000:00011:00001",
  "USGS:04119000:00011:00002",
  "USGS:04119055:00011:00002",
  "USGS:04119055:00011:00001",
  "USGS:04119400:00011:00006",
  "USGS:04119400:00011:00004",
  "USGS:04119400:00011:00002",
  "USGS:04119400:00011:00003",
  "USGS:04119400:00011:00007",
  "USGS:04119400:00011:00011",
  "USGS:04119400:00011:00008",
  "USGS:04119400:00011:00009",
  "USGS:04121300:00011:00001",
  "USGS:04121300:00011:00002",
  "USGS:04121500:00011:00001",
  "USGS:04121500:00011:00004",
  "USGS:04121650:00011:00003",
  "USGS:04121650:00011:00002",
  "USGS:04121660:00011:00001",
  "USGS:04121660:00011:00002",
  "USGS:04121680:00011:00001",
  "USGS:04121680:00011:00002",
  "USGS:04121944:00011:00005",
  "USGS:04121944:00011:00002",
  "USGS:04121944:00011:00001",
  "USGS:04121944:00011:00003",
  "USGS:04121970:00011:00003",
  "USGS:04121970:00011:00012",
  "USGS:04121970:00011:00001",
  "USGS:04121970:00011:00002",
  "USGS:04121970:00011:00008",
  "USGS:04121970:00011:00005",
  "USGS:04121970:00011:00009",
  "USGS:04121970:00011:00010",
  "USGS:04122100:00011:00001",
  "USGS:04122100:00011:00002",
  "USGS:04122200:00011:00001",
  "USGS:04122200:00011:00002",
  "USGS:0412220999:00011:00003",
  "USGS:0412220999:00011:00001",
  "USGS:0412220999:00011:00002",
  "USGS:04122500:00011:00001",
  "USGS:04122500:00011:00003",
  "USGS:04124000:00011:00003",
  "USGS:04124000:00011:00001",
  "USGS:04124000:00011:00002",
  "USGS:04124000:00011:00005",
  "USGS:04124200:00011:00003",
  "USGS:04124200:00011:00002",
  "USGS:04124200:00011:00001",
  "USGS:04124200:00011:00005",
  "USGS:04124500:00011:00001",
  "USGS:04124500:00011:00003",
  "USGS:04125460:00011:00003",
  "USGS:04125460:00011:00002",
  "USGS:04125460:00011:00001",
  "USGS:04125460:00011:00005",
  "USGS:04125550:00011:00004",
  "USGS:04125550:00011:00003",
  "USGS:04125550:00011:00002",
  "USGS:04125550:00011:00006",
  "USGS:04126740:00011:00002",
  "USGS:04126740:00011:00001",
  "USGS:04126970:00011:00003",
  "USGS:04126970:00011:00002",
  "USGS:04127800:00011:00001",
  "USGS:04127800:00011:00002",
  "USGS:04127885:00011:00004",
  "USGS:04127885:00011:00019",
  "USGS:04127917:00011:00001",
  "USGS:04127917:00011:00002",
  "USGS:04127997:00011:00002",
  "USGS:04127997:00011:00001",
  "USGS:04128990:00011:00002",
  "USGS:04128990:00011:00001",
  "USGS:04133501:00011:00002",
  "USGS:04133501:00011:00001",
  "USGS:04135700:00011:00002",
  "USGS:04135700:00011:00005",
  "USGS:04136000:00011:00004",
  "USGS:04136000:00011:00001",
  "USGS:04136000:00011:00008",
  "USGS:04136000:00011:00006",
  "USGS:05014300:00011:00003",
  "USGS:05014300:00011:00002",
  "USGS:05014300:00011:00001",
  "USGS:05014500:00011:00002",
  "USGS:05014500:00011:00006",
  "USGS:05015500:00011:00002",
  "USGS:05017500:00011:00001",
  "USGS:05017500:00011:00003",
  "USGS:05018000:00011:00001",
  "USGS:05018000:00011:00002",
  "USGS:05018500:00011:00001",
  "USGS:05018500:00011:00002",
  "USGS:01163200:00011:00001",
  "USGS:01163200:00011:00002",
  "USGS:01163500:00011:00003",
  "USGS:01163500:00011:00012",
  "USGS:01163500:00011:00001",
  "USGS:01163500:00011:00011",
  "USGS:01164000:00011:00001",
  "USGS:01164000:00011:00002",
  "USGS:01164000:00011:00011",
  "USGS:01165000:00011:00001",
  "USGS:01165000:00011:00008",
  "USGS:01166500:00011:00001",
  "USGS:01166500:00011:00005",
  "USGS:01168250:00011:00002",
  "USGS:01168500:00011:00001",
  "USGS:01168500:00011:00009",
  "USGS:01169000:00011:00001",
  "USGS:01169000:00011:00003",
  "USGS:01169900:00011:00001",
  "USGS:01169900:00011:00002",
  "USGS:01170000:00011:00007",
  "USGS:01170000:00011:00008",
  "USGS:01170100:00011:00015",
  "USGS:01170100:00011:00001",
  "USGS:01170100:00011:00003",
  "USGS:01170500:00011:00001",
  "USGS:01170500:00011:00005",
  "USGS:01171500:00011:00001",
  "USGS:01171500:00011:00002",
  "USGS:01172010:00011:00001",
  "USGS:01172010:00011:00002",
  "USGS:01172500:00011:00001",
  "USGS:01172500:00011:00005",
  "USGS:01173000:00011:00007",
  "USGS:01173000:00011:00001",
  "USGS:01173000:00011:00009",
  "USGS:01173500:00011:00001",
  "USGS:01173500:00011:00004",
  "USGS:01174500:00011:00001",
  "USGS:01174500:00011:00004",
  "USGS:01174565:00011:00001",
  "USGS:01174565:00011:00002",
  "USGS:01175500:00011:00013",
  "USGS:01175500:00011:00001",
  "USGS:01175500:00011:00002",
  "USGS:01175670:00011:00001",
  "USGS:01175670:00011:00002",
  "USGS:01176000:00011:00018",
  "USGS:01176000:00011:00001",
  "USGS:01176000:00011:00003",
  "USGS:01177000:00011:00001",
  "USGS:01177000:00011:00003",
  "USGS:01179500:00011:00001",
  "USGS:01179500:00011:00005",
  "USGS:01179500:00011:00008",
  "USGS:01180500:00011:00001",
  "USGS:01180500:00011:00005",
  "USGS:01181000:00011:00001",
  "USGS:01181000:00011:00003",
  "USGS:01183500:00011:00001",
  "USGS:01183500:00011:00004",
  "USGS:01185500:00011:00001",
  "USGS:01185500:00011:00006",
  "USGS:01197000:00011:00001",
  "USGS:01197000:00011:00003",
  "USGS:01197500:00011:00001",
  "USGS:01197500:00011:00005",
  "USGS:01198000:00011:00001",
  "USGS:01198000:00011:00002",
  "USGS:01198125:00011:00002",
  "USGS:01198125:00011:00001",
  "USGS:01331500:00011:00001",
  "USGS:01331500:00011:00002",
  "USGS:01332500:00011:00001",
  "USGS:01332500:00011:00004",
  "USGS:01333000:00011:00001",
  "USGS:01333000:00011:00002",
  "USGS:04015330:00011:00005",
  "USGS:04015330:00011:00004",
  "USGS:04015330:00011:00008",
  "USGS:04015330:00011:00006",
  "USGS:04015330:00011:00001",
  "USGS:04015330:00011:00009",
  "USGS:293229091230800:00011:00002",
  "USGS:293229091230800:00011:00001",
  "USGS:293229091230800:00011:00003",
  "USGS:293229091230800:00011:00005",
  "USGS:293229091230800:00011:00004",
  "USGS:413601070275800:00011:00002",
  "USGS:413601070275800:00011:00006",
  "USGS:413601070275800:00011:00004",
  "USGS:413601070275800:00011:00003",
  "USGS:413601070275800:00011:00007",
  "USGS:413601070275800:00011:00005",
  "USGS:413601070275800:00011:00001",
  "USGS:413758070320501:00011:00001",
  "USGS:05500000:00011:00007",
  "USGS:05500000:00011:00002",
  "USGS:05501000:00011:00003",
  "USGS:05501000:00011:00007",
  "USGS:05501000:00011:00002",
  "USGS:05501600:00011:00002",
  "USGS:05502000:00011:00001",
  "USGS:05502000:00011:00005",
  "USGS:05502300:00011:00003",
  "USGS:05502300:00011:00005",
  "USGS:05502300:00011:00002",
  "USGS:05502500:00011:00001",
  "USGS:05502500:00011:00003",
  "USGS:05503100:00011:00002",
  "USGS:05503100:00011:00001",
  "USGS:05503800:00011:00003",
  "USGS:05503800:00011:00005",
  "USGS:05503800:00011:00002",
  "USGS:05504800:00011:00001",
  "USGS:05504800:00011:00003",
  "USGS:05506100:00011:00012",
  "USGS:05506100:00011:00016",
  "USGS:05506100:00011:00001",
  "USGS:02475500:00011:00006",
  "USGS:07374000:00011:00015",
  "USGS:07374000:00011:00025",
  "USGS:07374000:00011:00020",
  "USGS:07374000:00011:00016",
  "USGS:07374000:00011:00028",
  "USGS:07374000:00011:00021",
  "USGS:07374000:00011:00031",
  "USGS:07374370:00011:00001",
  "USGS:07374510:00011:00001",
  "USGS:07374525:00011:00006",
  "USGS:07374525:00011:00019",
  "USGS:07374525:00011:00005",
  "USGS:07374525:00011:00023",
  "USGS:07374525:00011:00024",
  "USGS:073745253:00011:00001",
  "USGS:073745253:00011:00004",
  "USGS:073745253:00011:00002",
  "USGS:073745253:00011:00016",
  "USGS:073745253:00011:00017",
  "USGS:073745257:00011:00001",
  "USGS:073745257:00011:00004",
  "USGS:073745257:00011:00002",
  "USGS:073745257:00011:00014",
  "USGS:073745258:00011:00001",
  "USGS:073745258:00011:00004",
  "USGS:073745258:00011:00002",
  "USGS:073745258:00011:00014",
  "USGS:07374526:00011:00013",
  "USGS:07374526:00011:00001",
  "USGS:07374526:00011:00002",
  "USGS:07374526:00011:00014",
  "USGS:07374526:00011:00015",
  "USGS:07374527:00011:00015",
  "USGS:07374527:00011:00005",
  "USGS:07374527:00011:00006",
  "USGS:07374527:00011:00001",
  "USGS:07374527:00011:00002",
  "USGS:07374527:00011:00016",
  "USGS:07374527:00011:00018",
  "USGS:073745275:00011:00002",
  "USGS:073745275:00011:00001",
  "USGS:073745275:00011:00003",
  "USGS:073745275:00011:00004",
  "USGS:07374540:00011:00001",
  "USGS:07374540:00011:00002",
  "USGS:07374540:00011:00003",
  "USGS:07374550:00011:00001",
  "USGS:07374581:00011:00001",
  "USGS:07375000:00011:00001",
  "USGS:07375000:00011:00003",
  "USGS:07375000:00011:00015",
  "USGS:07375050:00011:00005",
  "USGS:07375050:00011:00004",
  "USGS:07375105:00011:00002",
  "USGS:07375105:00011:00001",
  "USGS:07375105:00011:00012",
  "USGS:07375175:00011:00002",
  "USGS:07375175:00011:00001",
  "USGS:07375175:00011:00012",
  "USGS:07375300:00011:00002",
  "USGS:07375300:00011:00001",
  "USGS:07375300:00011:00012",
  "USGS:07375430:00011:00002",
  "USGS:07375430:00011:00001",
  "USGS:07375430:00011:00012",
  "USGS:07375500:00011:00018",
  "USGS:07375500:00011:00019",
  "USGS:07375500:00011:00002",
  "USGS:07375500:00011:00005",
  "USGS:07375500:00011:00001",
  "USGS:07375500:00011:00022",
  "USGS:07375650:00011:00001",
  "USGS:07375800:00011:00014",
  "USGS:07375800:00011:00015",
  "USGS:07375800:00011:00002",
  "USGS:07375800:00011:00004",
  "USGS:07375800:00011:00001",
  "USGS:07375800:00011:00016",
  "USGS:07375960:00011:00002",
  "USGS:07375960:00011:00001",
  "USGS:07375960:00011:00012",
  "USGS:07376000:00011:00016",
  "USGS:07376000:00011:00017",
  "USGS:07376000:00011:00004",
  "USGS:07376000:00011:00001",
  "USGS:07376000:00011:00020",
  "USGS:07376500:00011:00005",
  "USGS:07376500:00011:00001",
  "USGS:07376500:00011:00004",
  "USGS:07376500:00011:00015",
  "USGS:07377000:00011:00004",
  "USGS:07377000:00011:00001",
  "USGS:07377000:00011:00019",
  "USGS:07377150:00011:00002",
  "USGS:07377150:00011:00001",
  "USGS:07377150:00011:00014",
  "USGS:07377195:00011:00001",
  "USGS:07377230:00011:00004",
  "USGS:07377230:00011:00003",
  "USGS:07377230:00011:00001",
  "USGS:07377300:00011:00001",
  "USGS:07377500:00011:00004",
  "USGS:07377500:00011:00002",
  "USGS:07377500:00011:00003",
  "USGS:07377500:00011:00018",
  "USGS:07377600:00011:00002",
  "USGS:07377600:00011:00001",
  "USGS:07377600:00011:00014",
  "USGS:07377750:00011:00002",
  "USGS:07377750:00011:00001",
  "USGS:07377750:00011:00014",
  "USGS:07377754:00011:00002",
  "USGS:07377754:00011:00001",
  "USGS:07377754:00011:00014",
  "USGS:07377760:00011:00002",
  "USGS:07377760:00011:00001",
  "USGS:07377760:00011:00012",
  "USGS:07377780:00011:00004",
  "USGS:07377780:00011:00003",
  "USGS:07377780:00011:00001",
  "USGS:07377870:00011:00002",
  "USGS:07377870:00011:00001",
  "USGS:07377870:00011:00014",
  "USGS:07378000:00011:00015",
  "USGS:07378000:00011:00014",
  "USGS:07378000:00011:00013",
  "USGS:07378000:00011:00020",
  "USGS:07378050:00011:00001",
  "USGS:07378083:00011:00002",
  "USGS:07378100:00011:00004",
  "USGS:07378100:00011:00003",
  "USGS:07378100:00011:00001",
  "USGS:293809092361500:00011:00002",
  "USGS:293809092361500:00011:00001",
  "USGS:293809092361500:00011:00003",
  "USGS:293809092361500:00011:00005",
  "USGS:293809092361500:00011:00004",
  "USGS:293809092361500:00011:00006",
  "USGS:06893791:00011:00017",
  "USGS:06893820:00011:00003",
  "USGS:06893820:00011:00005",
  "USGS:06893820:00011:00004",
  "USGS:06893820:00011:00002",
  "USGS:06893820:00011:00001",
  "USGS:06893820:00011:00006",
  "USGS:06893820:00011:00009",
  "USGS:06893820:00011:00008",
  "USGS:06893820:00011:00007",
  "USGS:06893820:00011:00010",
  "USGS:06893830:00011:00013",
  "USGS:07381600:00011:00023",
  "USGS:07381600:00011:00024",
  "USGS:07381600:00011:00001",
  "USGS:073816202:00011:00002",
  "USGS:073816501:00011:00001",
  "USGS:073816501:00011:00014",
  "USGS:073816503:00011:00002",
  "USGS:073816503:00011:00013",
  "USGS:073816503:00011:00015",
  "USGS:073816503:00011:00016",
  "USGS:07381670:00011:00002",
  "USGS:07381670:00011:00013",
  "USGS:07381670:00011:00001",
  "USGS:07382000:00011:00003",
  "USGS:07382000:00011:00006",
  "USGS:07382000:00011:00017",
  "USGS:07382500:00011:00018",
  "USGS:07382500:00011:00019",
  "USGS:07383500:00011:00002",
  "USGS:07383500:00011:00006",
  "USGS:07383500:00011:00017",
  "USGS:07383510:00011:00001",
  "USGS:07384400:00011:00002",
  "USGS:07385765:00011:00003",
  "USGS:07385765:00011:00004",
  "USGS:07385790:00011:00016",
  "USGS:07385790:00011:00014",
  "USGS:07385790:00011:00003",
  "USGS:07385820:00011:00001",
  "USGS:07386600:00011:00002",
  "USGS:07386600:00011:00001",
  "USGS:07386600:00011:00014",
  "USGS:07386850:00011:00001",
  "USGS:07386850:00011:00014",
  "USGS:07386880:00011:00020",
  "USGS:07386880:00011:00021",
  "USGS:07386880:00011:00017",
  "USGS:07386880:00011:00005",
  "USGS:07386880:00011:00014",
  "USGS:07386880:00011:00004",
  "USGS:07386880:00011:00019",
  "USGS:07386940:00011:00013",
  "USGS:07386940:00011:00001",
  "USGS:07386940:00011:00014",
  "USGS:07386980:00011:00001",
  "USGS:07386980:00011:00004",
  "USGS:07386980:00011:00006",
  "USGS:07386980:00011:00019",
  "USGS:07387040:00011:00006",
  "USGS:07387040:00011:00009",
  "USGS:07387040:00011:00010",
  "USGS:07387040:00011:00005",
  "USGS:07387040:00011:00007",
  "USGS:07387040:00011:00021",
  "USGS:07387040:00011:00028",
  "USGS:07387050:00011:00002",
  "USGS:07387050:00011:00001",
  "USGS:07387050:00011:00003",
  "USGS:07387050:00011:00016",
  "USGS:08010000:00011:00001",
  "USGS:08010000:00011:00003",
  "USGS:08012000:00011:00013",
  "USGS:08012000:00011:00014",
  "USGS:08012000:00011:00015",
  "USGS:08012000:00011:00001",
  "USGS:08012000:00011:00003",
  "USGS:08012000:00011:00016",
  "USGS:08012150:00011:00021",
  "USGS:08012150:00011:00018",
  "USGS:08012150:00011:00017",
  "USGS:08012150:00011:00022",
  "USGS:08013000:00011:00001",
  "USGS:08013000:00011:00003",
  "USGS:08013000:00011:00016",
  "USGS:08013500:00011:00003",
  "USGS:08013500:00011:00002",
  "USGS:08013500:00011:00001",
  "USGS:08013500:00011:00024",
  "USGS:08014500:00011:00017",
  "USGS:08014500:00011:00018",
  "USGS:08014500:00011:00019",
  "USGS:08014500:00011:00006",
  "USGS:08014500:00011:00001",
  "USGS:08014500:00011:00004",
  "USGS:08014500:00011:00020",
  "USGS:08014800:00011:00001",
  "USGS:08014800:00011:00002",
  "USGS:08014800:00011:00013",
  "USGS:08014881:00011:00001",
  "USGS:08014881:00011:00012",
  "USGS:08015500:00011:00019",
  "USGS:08015500:00011:00020",
  "USGS:08015500:00011:00008",
  "USGS:08015500:00011:00002",
  "USGS:08015500:00011:00006",
  "USGS:08017044:00011:00005",
  "USGS:08017044:00011:00003",
  "USGS:08017044:00011:00006",
  "USGS:08017044:00011:00024",
  "USGS:08017095:00011:00005",
  "USGS:08017095:00011:00008",
  "USGS:08017095:00011:00006",
  "USGS:08017095:00011:00018",
  "USGS:08017118:00011:00001",
  "USGS:08017118:00011:00005",
  "USGS:08017118:00011:00006",
  "USGS:08017118:00011:00004",
  "USGS:08017118:00011:00002",
  "USGS:08017118:00011:00017",
  "USGS:08023080:00011:00002",
  "USGS:08023080:00011:00007",
  "USGS:08023400:00011:00002",
  "USGS:08023400:00011:00007",
  "USGS:08025350:00011:00004",
  "USGS:08025350:00011:00001",
  "USGS:08025350:00011:00002",
  "USGS:08025500:00011:00001",
  "USGS:08025500:00011:00018",
  "USGS:08028000:00011:00002",
  "USGS:08028000:00011:00006",
  "USGS:291929089562600:00011:00004",
  "USGS:291929089562600:00011:00002",
  "USGS:291929089562600:00011:00015",
  "USGS:291929089562600:00011:00016",
  "USGS:292800090060000:00011:00002",
  "USGS:292800090060000:00011:00015",
  "USGS:292800090060000:00011:00016",
  "USGS:292800090060000:00011:00001",
  "USGS:292800090060000:00011:00003",
  "USGS:292800090060000:00011:00017",
  "USGS:292800090060000:00011:00018",
  "USGS:06917560:00011:00003",
  "USGS:06917560:00011:00002",
  "USGS:06917560:00011:00001",
  "USGS:06917630:00011:00005",
  "USGS:06917630:00011:00003",
  "USGS:06917630:00011:00002",
  "USGS:06917630:00011:00004",
  "USGS:06917630:00011:00006",
  "USGS:06917630:00011:00009",
  "USGS:06917630:00011:00007",
  "USGS:06918060:00011:00002",
  "USGS:06918060:00011:00001",
  "USGS:06918070:00011:00003",
  "USGS:06918250:00011:00018",
  "USGS:06918250:00011:00002",
  "USGS:06918250:00011:00001",
  "USGS:06918440:00011:00006",
  "USGS:06918440:00011:00002",
  "USGS:05355038:00011:00001",
  "USGS:05355080:00011:00001",
  "USGS:05355200:00011:00004",
  "USGS:05355200:00011:00003",
  "USGS:05372995:00011:00018",
  "USGS:05372995:00011:00007",
  "USGS:05372995:00011:00006",
  "USGS:05374000:00011:00003",
  "USGS:05378500:00011:00010",
  "USGS:05383950:00011:00002",
  "USGS:05383950:00011:00001",
  "USGS:05385000:00011:00008",
  "USGS:05385000:00011:00007",
  "USGS:05385500:00011:00002",
  "USGS:05385500:00011:00007",
  "USGS:05386400:00011:00001",
  "USGS:05457000:00011:00010",
  "USGS:05457000:00011:00014",
  "USGS:05475350:00011:00001",
  "USGS:05476000:00011:00002",
  "USGS:05476000:00011:00012",
  "USGS:05495000:00011:00003",
  "USGS:05495000:00011:00007",
  "USGS:05495000:00011:00002",
  "USGS:05496000:00011:00007",
  "USGS:05496000:00011:00002",
  "USGS:05497150:00011:00002",
  "USGS:05497150:00011:00001",
  "USGS:05498150:00011:00003",
  "USGS:05498150:00011:00002",
  "USGS:05498150:00011:00001",
  "USGS:05498700:00011:00012",
  "USGS:05498700:00011:00002",
  "USGS:05498700:00011:00001",
  "USGS:442917095183701:00011:00003",
  "USGS:442917095183701:00011:00006",
  "USGS:442917095183701:00011:00002",
  "USGS:442917095183701:00011:00001",
  "USGS:443912092423501:00011:00003",
  "USGS:443912092423501:00011:00001",
  "USGS:443912092423501:00011:00002",
  "USGS:443920092412701:00011:00002",
  "USGS:443920092412701:00011:00005",
  "USGS:443920092412701:00011:00008",
  "USGS:443920092412701:00011:00007",
  "USGS:443920092412702:00011:00002",
  "USGS:443920092412702:00011:00005",
  "USGS:443920092412702:00011:00004",
  "USGS:443920092412703:00011:00002",
  "USGS:443920092412703:00011:00005",
  "USGS:443920092412703:00011:00004",
  "USGS:444424095312301:00011:00002",
  "USGS:444424095312301:00011:00008",
  "USGS:444424095312301:00011:00007",
  "USGS:444431095324101:00011:00002",
  "USGS:444431095324101:00011:00005",
  "USGS:444431095324101:00011:00008",
  "USGS:444431095324101:00011:00007",
  "USGS:444443095305001:00011:00002",
  "USGS:444443095305001:00011:00008",
  "USGS:444443095305001:00011:00007",
  "USGS:444447095293501:00011:00002",
  "USGS:444447095293501:00011:00005",
  "USGS:444447095293501:00011:00004",
  "USGS:444447095293501:00011:00008",
  "USGS:444447095293501:00011:00007",
  "USGS:455927095123101:00011:00003",
  "USGS:455927095123101:00011:00005",
  "USGS:455927095123101:00011:00002",
  "USGS:455927095123101:00011:00001",
  "USGS:464646092052900:00011:00003",
  "USGS:464646092052900:00011:00001",
  "USGS:473423095053301:00011:00002",
  "USGS:473423095053301:00011:00006",
  "USGS:473423095053301:00011:00003",
  "USGS:473423095053301:00011:00001",
  "USGS:473841096153101:00011:00002",
  "USGS:473841096153101:00011:00005",
  "USGS:473841096153101:00011:00001",
  "USGS:473841096153101:00011:00006",
  "USGS:473933096243701:00011:00002",
  "USGS:473933096243701:00011:00005",
  "USGS:473933096243701:00011:00001",
  "USGS:473933096243701:00011:00006",
  "USGS:473945096202401:00011:00002",
  "USGS:473945096202401:00011:00001",
  "USGS:473945096202401:00011:00003",
  "USGS:473945096202402:00011:00002",
  "USGS:473945096202402:00011:00005",
  "USGS:473945096202402:00011:00001",
  "USGS:473945096202402:00011:00006",
  "USGS:474125096120602:00011:00002",
  "USGS:474125096120602:00011:00005",
  "USGS:474125096120602:00011:00001",
  "USGS:474125096120602:00011:00006",
  "USGS:474126096165301:00011:00002",
  "USGS:474126096165301:00011:00005",
  "USGS:474126096165301:00011:00001",
  "USGS:474126096165301:00011:00006",
  "USGS:474135096203001:00011:00002",
  "USGS:474135096203001:00011:00005",
  "USGS:474135096203001:00011:00001",
  "USGS:474135096203001:00011:00006",
  "USGS:474309096122001:00011:   NA",
  "USGS:474309096122001:00011:   NA",
  "USGS:474309096122001:00011:   NA",
  "USGS:474310096121801:00011:00002",
  "USGS:292952089453800:00011:00005",
  "USGS:474310096121801:00011:00005",
  "USGS:474310096121801:00011:00001",
  "USGS:474310096121801:00011:00006",
  "USGS:474346096185501:00011:00002",
  "USGS:474346096185501:00011:00005",
  "USGS:474346096185501:00011:00001",
  "USGS:474346096185501:00011:00006",
  "USGS:474436096140801:00011:00002",
  "USGS:474436096140801:00011:00008",
  "USGS:474436096140801:00011:00005",
  "USGS:474436096140801:00011:00001",
  "USGS:474436096140801:00011:00006",
  "USGS:474719096163100:00011:00002",
  "USGS:474719096163100:00011:00005",
  "USGS:474719096163100:00011:00001",
  "USGS:474719096163100:00011:00006",
  "USGS:474921093144001:00011:00012",
  "USGS:474921093144001:00011:00015",
  "USGS:474921093144001:00011:00011",
  "USGS:474921093144001:00011:00001",
  "USGS:06935755:00011:00002",
  "USGS:06935755:00011:00004",
  "USGS:06935770:00011:00003",
  "USGS:06935770:00011:00002",
  "USGS:06935830:00011:00002",
  "USGS:06935830:00011:00001",
  "USGS:06006000:00011:00002",
  "USGS:06006000:00011:00004",
  "USGS:06012500:00011:00005",
  "USGS:06012500:00011:00002",
  "USGS:06016000:00011:00002",
  "USGS:06016000:00011:00005",
  "USGS:06017000:00011:00001",
  "USGS:06017000:00011:00002",
  "USGS:06018500:00011:00005",
  "USGS:06018500:00011:00002",
  "USGS:06019500:00011:00001",
  "USGS:06019500:00011:00003",
  "USGS:06020600:00011:00001",
  "USGS:06020600:00011:00003",
  "USGS:06023000:00011:00001",
  "USGS:06023000:00011:00004",
  "USGS:06023000:00011:00005",
  "USGS:06023100:00011:00003",
  "USGS:06023100:00011:00002",
  "USGS:06023100:00011:00001",
  "USGS:06928380:00011:00002",
  "USGS:06928380:00011:00001",
  "USGS:292859090004000:00011:00002",
  "USGS:292859090004000:00011:00014",
  "USGS:292859090004000:00011:00003",
  "USGS:292859090004000:00011:00015",
  "USGS:292859090004000:00011:00016",
  "USGS:292952089453800:00011:00002",
  "USGS:292952089453800:00011:00001",
  "USGS:292952089453800:00011:00003",
  "USGS:292952089453800:00011:00004",
  "USGS:292952089453800:00011:00006",
  "USGS:292952090565300:00011:00002",
  "USGS:292952090565300:00011:00001",
  "USGS:292952090565300:00011:00003",
  "USGS:292952090565300:00011:00005",
  "USGS:292952090565300:00011:00004",
  "USGS:294736091164200:00011:00001",
  "USGS:295011091184300:00011:00002",
  "USGS:295011091184300:00011:00001",
  "USGS:2951190901217:00011:00002",
  "USGS:2951190901217:00011:00003",
  "USGS:2951190901217:00011:00015",
  "USGS:2951190901217:00011:00014",
  "USGS:295124089542100:00011:00012",
  "USGS:295124089542100:00011:00002",
  "USGS:295124089542100:00011:00013",
  "USGS:295124089542100:00011:00001",
  "USGS:295124089542100:00011:00014",
  "USGS:295124089542100:00011:00016",
  "USGS:295124089542100:00011:00017",
  "USGS:295231093100100:00011:00002",
  "USGS:295231093100100:00011:00001",
  "USGS:295231093100100:00011:00003",
  "USGS:295231093100100:00011:00005",
  "USGS:295231093100100:00011:00004",
  "USGS:295231093100100:00011:00006",
  "USGS:295447091191500:00011:00002",
  "USGS:295447091191500:00011:00001",
  "USGS:295501090190400:00011:00003",
  "USGS:295501090190400:00011:00002",
  "USGS:295501090190400:00011:00017",
  "USGS:295501090190400:00011:00001",
  "USGS:295501090190400:00011:00004",
  "USGS:295501090190400:00011:00016",
  "USGS:295501090190400:00011:00015",
  "USGS:295744093303800:00011:00002",
  "USGS:295744093303800:00011:00001",
  "USGS:295744093303800:00011:00003",
  "USGS:295744093303800:00011:00005",
  "USGS:295744093303800:00011:00004",
  "USGS:295744093303800:00011:00006",
  "USGS:295827090052800:00011:00002",
  "USGS:295827090052800:00011:00001",
  "USGS:295827090052800:00011:00003",
  "USGS:295827090052800:00011:00007",
  "USGS:295827090052800:00011:00005",
  "USGS:295827090052800:00011:00004",
  "USGS:295827090052800:00011:00006",
  "USGS:295906090054200:00011:00002",
  "USGS:295906090054200:00011:00001",
  "USGS:295906090054200:00011:00003",
  "USGS:295906090054200:00011:00007",
  "USGS:295906090054200:00011:00005",
  "USGS:295906090054200:00011:00004",
  "USGS:295906090054200:00011:00006",
  "USGS:300009090051600:00011:00002",
  "USGS:300009090051600:00011:00001",
  "USGS:300009090051600:00011:00003",
  "USGS:300009090051600:00011:00007",
  "USGS:300009090051600:00011:00005",
  "USGS:300009090051600:00011:00004",
  "USGS:300009090051600:00011:00006",
  "USGS:300026090050800:00011:00002",
  "USGS:300026090050800:00011:00001",
  "USGS:300026090050800:00011:00003",
  "USGS:300026090050800:00011:00007",
  "USGS:300026090050800:00011:00005",
  "USGS:300026090050800:00011:00004",
  "USGS:300026090050800:00011:00006",
  "USGS:300034090055300:00011:00002",
  "USGS:300034090055300:00011:00012",
  "USGS:300034090055300:00011:00014",
  "USGS:300034090055300:00011:00009",
  "USGS:300034090055300:00011:00010",
  "USGS:300034090055300:00011:00011",
  "USGS:300034090055300:00011:00008",
  "USGS:300034090055300:00011:00013",
  "USGS:300034090055300:00011:00001",
  "USGS:300034090055300:00011:00003",
  "USGS:300034090055300:00011:00007",
  "USGS:300034090055300:00011:00005",
  "USGS:300034090055300:00011:00004",
  "USGS:300034090055300:00011:00006",
  "USGS:300127090045800:00011:00002",
  "USGS:300127090045800:00011:00001",
  "USGS:300127090045800:00011:00003",
  "USGS:300127090045800:00011:00007",
  "USGS:300127090045800:00011:00005",
  "USGS:300127090045800:00011:00004",
  "USGS:300127090045800:00011:00006",
  "USGS:300128090045800:00011:00002",
  "USGS:300128090045800:00011:00001",
  "USGS:300128090045800:00011:00003",
  "USGS:300128090045800:00011:00007",
  "USGS:300128090045800:00011:00005",
  "USGS:300128090045800:00011:00004",
  "USGS:300128090045800:00011:00006",
  "USGS:300312091320000:00011:00002",
  "USGS:300312091320000:00011:00001",
  "USGS:300507091355600:00011:00003",
  "USGS:300507091355600:00011:00002",
  "USGS:300507091355600:00011:00001",
  "USGS:300602090375100:00011:00002",
  "USGS:300602090375100:00011:00001",
  "USGS:300602090375100:00011:00003",
  "USGS:300602090375100:00011:00005",
  "USGS:300602090375100:00011:00004",
  "USGS:300602090375100:00011:00006",
  "USGS:300713091362400:00011:00003",
  "USGS:300713091362400:00011:00002",
  "USGS:300713091362400:00011:00001",
  "USGS:300722089150100:00011:00001",
  "USGS:300722089150100:00011:00006",
  "USGS:300722089150100:00011:00005",
  "USGS:300722089150100:00011:00004",
  "USGS:300722089150100:00011:00002",
  "USGS:300722089150100:00011:00017",
  "USGS:301001089442600:00011:00003",
  "USGS:301001089442600:00011:00001",
  "USGS:301001089442600:00011:00004",
  "USGS:301001089442600:00011:00005",
  "USGS:301300092584503:00011:00001",
  "USGS:301324090382400:00011:00002",
  "USGS:301324090382400:00011:00001",
  "USGS:301324090382400:00011:00003",
  "USGS:301324090382400:00011:00005",
  "USGS:301324090382400:00011:00004",
  "USGS:301324090382400:00011:00006",
  "USGS:301655091440800:00011:00001",
  "USGS:301655091440800:00011:00012",
  "USGS:302020091435700:00011:00001",
  "USGS:302020091435700:00011:00012",
  "USGS:302614091083001:00011:00001",
  "USGS:302636091083802:00011:00001",
  "USGS:302642091083401:00011:00001",
  "USGS:321338092345801:00011:00001",
  "USGS:324141092390501:00011:00001",
  "USGS:330002092445901:00011:00001",
  "USGS:06079000:00011:00001",
  "USGS:06079000:00011:00002",
  "USGS:07019317:00011:00002",
  "USGS:07019317:00011:00001",
  "USGS:07020550:00011:00002",
  "USGS:07020550:00011:00001",
  "USGS:07020850:00011:00005",
  "USGS:05212700:00011:00002",
  "USGS:05227500:00011:00004",
  "USGS:05227500:00011:00003",
  "USGS:05227530:00011:00002",
  "USGS:05227530:00011:00001",
  "USGS:05242300:00011:00010",
  "USGS:05242300:00011:00009",
  "USGS:05243725:00011:00008",
  "USGS:05243725:00011:00007",
  "USGS:05244000:00011:00007",
  "USGS:05244000:00011:00003",
  "USGS:05245100:00011:00004",
  "USGS:05245100:00011:00006",
  "USGS:05247500:00011:00001",
  "USGS:05247500:00011:00007",
  "USGS:05267000:00011:00002",
  "USGS:05267000:00011:00007",
  "USGS:05270500:00011:00005",
  "USGS:05270500:00011:00004",
  "USGS:05270700:00011:00004",
  "USGS:05270700:00011:00003",
  "USGS:05275000:00011:00007",
  "USGS:05275000:00011:00002",
  "USGS:05280000:00011:00008",
  "USGS:05280000:00011:00007",
  "USGS:05280000:00011:00031",
  "USGS:05284000:00011:00005",
  "USGS:05286000:00011:00017",
  "USGS:05286000:00011:00001",
  "USGS:05287890:00011:00006",
  "USGS:05287890:00011:00003",
  "USGS:05288500:00011:00010",
  "USGS:05288500:00011:00006",
  "USGS:05288580:00011:00002",
  "USGS:05288580:00011:00001",
  "USGS:05288705:00011:00004",
  "USGS:05288705:00011:00002",
  "USGS:05288705:00011:00001",
  "USGS:05288705:00011:00005",
  "USGS:05289800:00011:00013",
  "USGS:05289800:00011:00003",
  "USGS:05289800:00011:00002",
  "USGS:05289800:00011:00001",
  "USGS:05289800:00011:00014",
  "USGS:05292000:00011:00004",
  "USGS:05292000:00011:00003",
  "USGS:05293000:00011:00019",
  "USGS:05293000:00011:00002",
  "USGS:05293000:00011:00007",
  "USGS:05294000:00011:00001",
  "USGS:05294000:00011:00004",
  "USGS:05294000:00011:00003",
  "USGS:05300000:00011:00004",
  "USGS:05300000:00011:00003",
  "USGS:05301000:00011:00005",
  "USGS:05301000:00011:00004",
  "USGS:05304500:00011:00008",
  "USGS:05304500:00011:00007",
  "USGS:05304995:00011:00001",
  "USGS:05305000:00011:00001",
  "USGS:05305000:00011:00003",
  "USGS:05311000:00011:00005",
  "USGS:05311000:00011:00004",
  "USGS:05311150:00011:00002",
  "USGS:05311150:00011:00001",
  "USGS:05313500:00011:00007",
  "USGS:05313500:00011:00009",
  "USGS:05315000:00011:00009",
  "USGS:05315000:00011:00020",
  "USGS:05316500:00011:00009",
  "USGS:05316500:00011:00012",
  "USGS:05316580:00011:00002",
  "USGS:05316580:00011:00001",
  "USGS:05317000:00011:00008",
  "USGS:05317000:00011:00007",
  "USGS:05317200:00011:00004",
  "USGS:05317200:00011:00003",
  "USGS:05319500:00011:00006",
  "USGS:05319500:00011:00007",
  "USGS:05320000:00011:00004",
  "USGS:05320000:00011:00003",
  "USGS:05320500:00011:00004",
  "USGS:05320500:00011:00002",
  "USGS:05325000:00011:00009",
  "USGS:05325000:00011:00014",
  "USGS:05325000:00011:00013",
  "USGS:05327000:00011:00004",
  "USGS:05327000:00011:00005",
  "USGS:05330000:00011:00007",
  "USGS:05330000:00011:00003",
  "USGS:05330000:00011:00006",
  "USGS:05330920:00011:00007",
  "USGS:05330920:00011:00021",
  "USGS:05330920:00011:00002",
  "USGS:05330920:00011:00006",
  "USGS:05331000:00011:00002",
  "USGS:05331000:00011:00004",
  "USGS:05331580:00011:   NA",
  "USGS:05331580:00011:   NA",
  "USGS:05331580:00011:   NA",
  "USGS:05331580:00011:   NA",
  "USGS:05336700:00011:00004",
  "USGS:05336700:00011:00003",
  "USGS:07068000:00011:00006",
  "USGS:07068000:00011:00002",
  "USGS:07068510:00011:00002",
  "USGS:07068510:00011:00003",
  "USGS:07071000:00011:00001",
  "USGS:07071000:00011:00007",
  "USGS:07071500:00011:00005",
  "USGS:07071500:00011:00002",
  "USGS:07185700:00011:00001",
  "USGS:07185700:00011:00002",
  "USGS:07185765:00011:00016",
  "USGS:07185765:00011:00001",
  "USGS:07185765:00011:00002",
  "USGS:07185910:00011:00002",
  "USGS:07185910:00011:00001",
  "USGS:07186000:00011:00005",
  "USGS:07186000:00011:00002",
  "USGS:07186480:00011:00002",
  "USGS:07186480:00011:00001",
  "USGS:07378500:00011:00009",
  "USGS:07378500:00011:00003",
  "USGS:07378500:00011:00005",
  "USGS:07378500:00011:00001",
  "USGS:07378500:00011:00020",
  "USGS:07378650:00011:00004",
  "USGS:07378650:00011:00003",
  "USGS:07378650:00011:00002",
  "USGS:07378722:00011:00004",
  "USGS:07378722:00011:00003",
  "USGS:07378722:00011:00014",
  "USGS:07378745:00011:00001",
  "USGS:07378745:00011:00003",
  "USGS:07378746:00011:00003",
  "USGS:07378746:00011:00001",
  "USGS:07378746:00011:00016",
  "USGS:07378748:00011:00001",
  "USGS:07378748:00011:00012",
  "USGS:07378810:00011:00004",
  "USGS:07378810:00011:00003",
  "USGS:07378810:00011:00014",
  "USGS:07379000:00011:00003",
  "USGS:07379050:00011:00005",
  "USGS:07379050:00011:00004",
  "USGS:07379050:00011:00015",
  "USGS:07379100:00011:00004",
  "USGS:07379100:00011:00003",
  "USGS:07379960:00011:00008",
  "USGS:07379960:00011:00007",
  "USGS:07379960:00011:00020",
  "USGS:07380101:00011:00002",
  "USGS:07380101:00011:00015",
  "USGS:07380102:00011:00004",
  "USGS:07380102:00011:00003",
  "USGS:07380102:00011:00015",
  "USGS:07380107:00011:00002",
  "USGS:07380107:00011:00001",
  "USGS:07380107:00011:00014",
  "USGS:073801175:00011:00001",
  "USGS:073801175:00011:00014",
  "USGS:07380120:00011:00018",
  "USGS:07380120:00011:00006",
  "USGS:07380120:00011:00015",
  "USGS:07380120:00011:00004",
  "USGS:07380120:00011:00025",
  "USGS:07380126:00011:00002",
  "USGS:07380126:00011:00001",
  "USGS:07380126:00011:00014",
  "USGS:07380144:00011:00001",
  "USGS:07380185:00011:00001",
  "USGS:07380185:00011:00014",
  "USGS:07380200:00011:00004",
  "USGS:07380200:00011:00003",
  "USGS:07380200:00011:00014",
  "USGS:07380215:00011:00003",
  "USGS:07380215:00011:00004",
  "USGS:07380215:00011:00002",
  "USGS:07380215:00011:00001",
  "USGS:07380215:00011:00014",
  "USGS:073802220:00011:00002",
  "USGS:073802220:00011:00001",
  "USGS:073802220:00011:00014",
  "USGS:073802225:00011:00003",
  "USGS:073802225:00011:00001",
  "USGS:073802225:00011:00002",
  "USGS:0738022295:00011:00002",
  "USGS:0738022295:00011:00001",
  "USGS:0738022295:00011:00015",
  "USGS:0738022395:00011:00002",
  "USGS:0738022395:00011:00001",
  "USGS:0738022395:00011:00014",
  "USGS:073802245:00011:00002",
  "USGS:073802245:00011:00001",
  "USGS:073802245:00011:00013",
  "USGS:073802273:00011:00002",
  "USGS:073802273:00011:00001",
  "USGS:073802273:00011:00013",
  "USGS:073802282:00011:00003",
  "USGS:073802282:00011:00001",
  "USGS:073802282:00011:00002",
  "USGS:073802332:00011:00002",
  "USGS:073802332:00011:00001",
  "USGS:07380238:00011:00002",
  "USGS:07380238:00011:00003",
  "USGS:07380238:00011:00013",
  "USGS:07380251:00011:00005",
  "USGS:07380251:00011:00010",
  "USGS:07380251:00011:00011",
  "USGS:07380251:00011:00008",
  "USGS:07380251:00011:00006",
  "USGS:07380251:00011:00021",
  "USGS:07380251:00011:00023",
  "USGS:073802512:00011:00006",
  "USGS:073802512:00011:00005",
  "USGS:073802512:00011:00007",
  "USGS:073802512:00011:00019",
  "USGS:073802512:00011:00020",
  "USGS:073802516:00011:00002",
  "USGS:073802516:00011:00005",
  "USGS:073802516:00011:00006",
  "USGS:073802516:00011:00001",
  "USGS:073802516:00011:00024",
  "USGS:073802516:00011:00003",
  "USGS:073802516:00011:00004",
  "USGS:073802516:00011:00021",
  "USGS:07380330:00011:00002",
  "USGS:07380330:00011:00001",
  "USGS:07380330:00011:00003",
  "USGS:07380330:00011:00004",
  "USGS:07380335:00011:00006",
  "USGS:07380335:00011:00005",
  "USGS:07380335:00011:00007",
  "USGS:07380335:00011:00019",
  "USGS:07380400:00011:00005",
  "USGS:07380400:00011:00006",
  "USGS:07380400:00011:00002",
  "USGS:07380401:00011:00014",
  "USGS:07352000:00011:00002",
  "USGS:07380401:00011:00012",
  "USGS:07380401:00011:00001",
  "USGS:07380401:00011:00015",
  "USGS:07380500:00011:00001",
  "USGS:07381000:00011:00015",
  "USGS:07381000:00011:00005",
  "USGS:07381000:00011:00003",
  "USGS:07381000:00011:00016",
  "USGS:07381150:00011:00002",
  "USGS:07381150:00011:00001",
  "USGS:07381150:00011:00003",
  "USGS:07381150:00011:00013",
  "USGS:07381150:00011:00014",
  "USGS:07381235:00011:00003",
  "USGS:07381235:00011:00002",
  "USGS:07381235:00011:00017",
  "USGS:07381235:00011:00001",
  "USGS:07381235:00011:00004",
  "USGS:07381235:00011:00016",
  "USGS:07381235:00011:00018",
  "USGS:07381324:00011:00019",
  "USGS:07381324:00011:00005",
  "USGS:07381324:00011:00015",
  "USGS:07381324:00011:00004",
  "USGS:07381324:00011:00017",
  "USGS:07381324:00011:00020",
  "USGS:07381324:00011:00021",
  "USGS:07381328:00011:00007",
  "USGS:07381328:00011:00016",
  "USGS:07381328:00011:00017",
  "USGS:07381328:00011:00009",
  "USGS:07381328:00011:00023",
  "USGS:07381328:00011:00018",
  "USGS:07381328:00011:00003",
  "USGS:07381328:00011:00001",
  "USGS:07381328:00011:00019",
  "USGS:07381328:00011:00021",
  "USGS:07381349:00011:00005",
  "USGS:07381349:00011:00009",
  "USGS:07381349:00011:00010",
  "USGS:07381349:00011:00008",
  "USGS:07381349:00011:00006",
  "USGS:07381349:00011:00018",
  "USGS:073813498:00011:00002",
  "USGS:073813498:00011:00005",
  "USGS:073813498:00011:00006",
  "USGS:073813498:00011:00001",
  "USGS:073813498:00011:00003",
  "USGS:073813498:00011:00019",
  "USGS:07381350:00011:00001",
  "USGS:07381350:00011:00003",
  "USGS:07381350:00011:00002",
  "USGS:07381350:00011:00014",
  "USGS:07381350:00011:00015",
  "USGS:07381355:00011:00002",
  "USGS:07381355:00011:00001",
  "USGS:07381355:00011:00003",
  "USGS:07381355:00011:00014",
  "USGS:07381355:00011:00015",
  "USGS:07381450:00011:00003",
  "USGS:07381454:00011:00001",
  "USGS:294045092492300:00011:00002",
  "USGS:294045092492300:00011:00001",
  "USGS:294045092492300:00011:00003",
  "USGS:294045092492300:00011:00005",
  "USGS:294045092492300:00011:00004",
  "USGS:294045092492300:00011:00006",
  "USGS:323830088491200:00011:00001",
  "USGS:370224094320201:00011:00001",
  "USGS:370236093174401:00011:00001",
  "USGS:370248090042601:00011:00002",
  "USGS:370354093325901:00011:00001",
  "USGS:370539093494001:00011:00011",
  "USGS:370539093494001:00011:00001",
  "USGS:370539093494002:00011:00001",
  "USGS:370600094223501:00011:00002",
  "USGS:370624092244701:00011:00011",
  "USGS:370624092244701:00011:00001",
  "USGS:370655093035301:00011:00001",
  "USGS:370828094274101:00011:00001",
  "USGS:370907093144101:00011:00001",
  "USGS:371036094171301:00011:00001",
  "USGS:371125089445301:00011:00002",
  "USGS:371220094302401:00011:00001",
  "USGS:371435093134701:00011:00001",
  "USGS:371548093144701:00011:00012",
  "USGS:371548093144701:00011:00001",
  "USGS:371548093144702:00011:00001",
  "USGS:371558093181901:00011:00001",
  "USGS:371800092094801:00011:00001",
  "USGS:07349298:00011:00012",
  "USGS:07349450:00011:00002",
  "USGS:07349500:00011:00004",
  "USGS:07349500:00011:00014",
  "USGS:07349650:00011:00001",
  "USGS:07349660:00011:00001",
  "USGS:07349815:00011:00001",
  "USGS:07349815:00011:00013",
  "USGS:07349849:00011:00001",
  "USGS:07349849:00011:00012",
  "USGS:07349860:00011:00001",
  "USGS:07349860:00011:00003",
  "USGS:07349860:00011:00014",
  "USGS:07349898:00011:00001",
  "USGS:07349898:00011:00012",
  "USGS:07349910:00011:00001",
  "USGS:07349910:00011:00012",
  "USGS:07350700:00011:00001",
  "USGS:07350700:00011:00013",
  "USGS:07350985:00011:00001",
  "USGS:07350985:00011:00013",
  "USGS:07351275:00011:00001",
  "USGS:07351275:00011:00012",
  "USGS:07351500:00011:00001",
  "USGS:07351500:00011:00003",
  "USGS:07351500:00011:00016",
  "USGS:07351550:00011:00001",
  "USGS:07351750:00011:00001",
  "USGS:07351750:00011:00007",
  "USGS:07351755:00011:00001",
  "USGS:07352000:00011:00006",
  "USGS:07352820:00011:00001",
  "USGS:07352820:00011:00002",
  "USGS:07352895:00011:00002",
  "USGS:07352895:00011:00013",
  "USGS:07353520:00011:00013",
  "USGS:07353520:00011:00001",
  "USGS:07364200:00011:00002",
  "USGS:07364200:00011:00008",
  "USGS:07364203:00011:00001",
  "USGS:07364300:00011:00002",
  "USGS:07364535:00011:00025",
  "USGS:07364840:00011:00014",
  "USGS:07364840:00011:00001",
  "USGS:07366200:00011:00002",
  "USGS:07366200:00011:00008",
  "USGS:07366364:00011:00012",
  "USGS:07366364:00011:00001",
  "USGS:07366472:00011:00003",
  "USGS:07367005:00011:00014",
  "USGS:07367005:00011:00003",
  "USGS:07367005:00011:00002",
  "USGS:07367005:00011:00001",
  "USGS:07367005:00011:00018",
  "USGS:07367690:00011:00002",
  "USGS:07367690:00011:00001",
  "USGS:07368000:00011:00002",
  "USGS:07368000:00011:00008",
  "USGS:07369000:00011:00005",
  "USGS:07369000:00011:00001",
  "USGS:07369050:00011:00004",
  "USGS:07369500:00011:00005",
  "USGS:07369500:00011:00001",
  "USGS:07369515:00011:00001",
  "USGS:375920092463001:00011:00001",
  "USGS:375930094222001:00011:00015",
  "USGS:375930094222001:00011:00013",
  "USGS:375930094222001:00011:00012",
  "USGS:375930094222001:00011:00011",
  "USGS:375930094222001:00011:00016",
  "USGS:375930094222001:00011:00014",
  "USGS:375930094222001:00011:00017",
  "USGS:375930094222001:00011:00019",
  "USGS:375930094222001:00011:00001",
  "USGS:380038092442701:00011:00001",
  "USGS:380229093464701:00011:00002",
  "USGS:380322091142601:00011:00001",
  "USGS:380435090281301:00011:00001",
  "USGS:380501090335501:00011:00002",
  "USGS:380545094213501:00011:00011",
  "USGS:380545094213501:00011:00001",
  "USGS:380717092395401:00011:00001",
  "USGS:380900091153901:00011:00001",
  "USGS:381045091564801:00011:00001",
  "USGS:381217091104501:00011:00001",
  "USGS:381405090260301:00011:00001",
  "USGS:381641093214601:00011:00011",
  "USGS:381641093214601:00011:00001",
  "USGS:381652093215501:00011:00002",
  "USGS:382100090592801:00011:00002",
  "USGS:06893830:00011:00014",
  "USGS:06893830:00011:00003",
  "USGS:06893830:00011:00002",
  "USGS:06893830:00011:00001",
  "USGS:06893830:00011:00016",
  "USGS:06893830:00011:00019",
  "USGS:06893885:00011:00015",
  "USGS:06893890:00011:00030",
  "USGS:06893890:00011:00016",
  "USGS:06893890:00011:00015",
  "USGS:06893890:00011:00001",
  "USGS:06893890:00011:00004",
  "USGS:06893890:00011:00018",
  "USGS:06893890:00011:00019",
  "USGS:06893890:00011:00031",
  "USGS:06893890:00011:00017",
  "USGS:06893890:00011:00020",
  "USGS:06893970:00011:00010",
  "USGS:06893970:00011:00004",
  "USGS:06893970:00011:00003",
  "USGS:06893970:00011:00002",
  "USGS:06893970:00011:00001",
  "USGS:06893970:00011:00006",
  "USGS:06893970:00011:00008",
  "USGS:06893970:00011:00009",
  "USGS:06893970:00011:00005",
  "USGS:06893970:00011:00007",
  "USGS:06894000:00011:00017",
  "USGS:06894000:00011:00016",
  "USGS:06894000:00011:00014",
  "USGS:06894000:00011:00004",
  "USGS:06894000:00011:00002",
  "USGS:06894000:00011:00019",
  "USGS:06894000:00011:00021",
  "USGS:06894000:00011:00022",
  "USGS:06894000:00011:00018",
  "USGS:06894000:00011:00020",
  "USGS:06894200:00011:00002",
  "USGS:06894200:00011:00001",
  "USGS:06894650:00011:00001",
  "USGS:06895000:00011:00001",
  "USGS:06895000:00011:00002",
  "USGS:06895500:00011:00005",
  "USGS:06895500:00011:00002",
  "USGS:06896000:00011:00012",
  "USGS:06896000:00011:00001",
  "USGS:06896000:00011:00002",
  "USGS:06896189:00011:00011",
  "USGS:06896189:00011:00012",
  "USGS:06896189:00011:00001",
  "USGS:06896400:00011:00003",
  "USGS:06896400:00011:00002",
  "USGS:06896400:00011:00001",
  "USGS:06896900:00011:00001",
  "USGS:06897000:00011:00016",
  "USGS:06897000:00011:00001",
  "USGS:06897000:00011:00003",
  "USGS:06897500:00011:00015",
  "USGS:06897500:00011:00004",
  "USGS:06897500:00011:00002",
  "USGS:06899500:00011:00004",
  "USGS:06899500:00011:00002",
  "USGS:06899680:00011:00002",
  "USGS:06899700:00011:00001",
  "USGS:06899700:00011:00002",
  "USGS:06899900:00011:00003",
  "USGS:06899900:00011:00002",
  "USGS:06899900:00011:00001",
  "USGS:06900050:00011:00013",
  "USGS:06900050:00011:00001",
  "USGS:06900640:00011:00004",
  "USGS:06900640:00011:00002",
  "USGS:06900640:00011:00001",
  "USGS:06901205:00011:00002",
  "USGS:06901205:00011:00001",
  "USGS:06901250:00011:00005",
  "USGS:06901250:00011:00003",
  "USGS:06901250:00011:00001",
  "USGS:06901500:00011:00016",
  "USGS:06901500:00011:00001",
  "USGS:06901500:00011:00002",
  "USGS:06902000:00011:00005",
  "USGS:06902000:00011:00002",
  "USGS:06902100:00011:00003",
  "USGS:06902990:00011:00011",
  "USGS:06902990:00011:00012",
  "USGS:06902990:00011:00001",
  "USGS:06902995:00011:00004",
  "USGS:06902995:00011:00002",
  "USGS:06902995:00011:00001",
  "USGS:06904050:00011:00003",
  "USGS:06904050:00011:00004",
  "USGS:06904050:00011:00002",
  "USGS:06904500:00011:00003",
  "USGS:06904500:00011:00005",
  "USGS:06904500:00011:00002",
  "USGS:06904500:00011:00018",
  "USGS:06905500:00011:00003",
  "USGS:06905500:00011:00006",
  "USGS:06905500:00011:00002",
  "USGS:06906000:00011:00015",
  "USGS:06906000:00011:00001",
  "USGS:06906000:00011:00003",
  "USGS:06906150:00011:00021",
  "USGS:06906150:00011:00001",
  "USGS:06906190:00011:00016",
  "USGS:06906200:00011:00001",
  "USGS:06906200:00011:00003",
  "USGS:06906500:00011:00019",
  "USGS:06906500:00011:00017",
  "USGS:06906500:00011:00002",
  "USGS:06906800:00011:00014",
  "USGS:06906800:00011:00002",
  "USGS:06906800:00011:00003",
  "USGS:06907700:00011:00003",
  "USGS:06907700:00011:00001",
  "USGS:06907700:00011:00002",
  "USGS:06907720:00011:00011",
  "USGS:06907720:00011:00012",
  "USGS:06907720:00011:00001",
  "USGS:06908000:00011:00004",
  "USGS:06908000:00011:00002",
  "USGS:06909000:00011:00006",
  "USGS:06909000:00011:00002",
  "USGS:06909500:00011:00015",
  "USGS:06909500:00011:00001",
  "USGS:06909500:00011:00002",
  "USGS:06909950:00011:00003",
  "USGS:06909950:00011:00002",
  "USGS:06909950:00011:00001",
  "USGS:06910230:00011:00002",
  "USGS:06910230:00011:00003",
  "USGS:06910450:00011:00012",
  "USGS:06910450:00011:00034",
  "USGS:06910450:00011:00001",
  "USGS:06910750:00011:00015",
  "USGS:06910750:00011:00001",
  "USGS:06910750:00011:00003",
  "USGS:06917060:00011:00013",
  "USGS:06917060:00011:00001",
  "USGS:10254730:00011:00007",
  "USGS:10254730:00011:00009",
  "USGS:10254730:00011:00001",
  "USGS:10254730:00011:00006",
  "USGS:02435020:00011:00008",
  "USGS:02436500:00011:00004",
  "USGS:02436500:00011:00003",
  "USGS:02437000:00011:00005",
  "USGS:02437000:00011:00004",
  "USGS:02437100:00011:00001",
  "USGS:06918460:00011:00005",
  "USGS:06918460:00011:00002",
  "USGS:06918493:00011:00024",
  "USGS:06918493:00011:00002",
  "USGS:06918493:00011:00003",
  "USGS:06918740:00011:00004",
  "USGS:06918740:00011:00002",
  "USGS:06918990:00011:00007",
  "USGS:06919000:00011:00003",
  "USGS:06919020:00011:00004",
  "USGS:06919020:00011:00002",
  "USGS:06919500:00011:00004",
  "USGS:06919500:00011:00002",
  "USGS:06919900:00011:00005",
  "USGS:06919900:00011:00002",
  "USGS:06920520:00011:00002",
  "USGS:06920520:00011:00001",
  "USGS:06921070:00011:00016",
  "USGS:06921070:00011:00005",
  "USGS:06921070:00011:00002",
  "USGS:06921200:00011:00005",
  "USGS:06921200:00011:00002",
  "USGS:06921325:00011:00010",
  "USGS:06921350:00011:00002",
  "USGS:06921350:00011:00017",
  "USGS:06921590:00011:00003",
  "USGS:06921590:00011:00005",
  "USGS:06921590:00011:00002",
  "USGS:06921600:00011:00002",
  "USGS:06921720:00011:00012",
  "USGS:06921720:00011:00001",
  "USGS:06921720:00011:00002",
  "USGS:06921760:00011:00005",
  "USGS:06921760:00011:00003",
  "USGS:06922440:00011:00003",
  "USGS:06922500:00011:00003",
  "USGS:06923250:00011:00002",
  "USGS:06923250:00011:00001",
  "USGS:06923500:00011:00002",
  "USGS:06923500:00011:00003",
  "USGS:06923940:00011:00002",
  "USGS:06923940:00011:00001",
  "USGS:06923950:00011:00016",
  "USGS:06923950:00011:00015",
  "USGS:06923950:00011:00001",
  "USGS:06925250:00011:00002",
  "USGS:06925250:00011:00001",
  "USGS:06926000:00011:00001",
  "USGS:06926000:00011:00003",
  "USGS:06926290:00011:00012",
  "USGS:06926290:00011:00002",
  "USGS:06926290:00011:00001",
  "USGS:06926510:00011:00016",
  "USGS:06926510:00011:00004",
  "USGS:06926510:00011:00005",
  "USGS:06927000:00011:00001",
  "USGS:06927000:00011:00002",
  "USGS:06927240:00011:00002",
  "USGS:06927240:00011:00001",
  "USGS:06928000:00011:00016",
  "USGS:06928000:00011:00001",
  "USGS:06928000:00011:00002",
  "USGS:06928300:00011:00016",
  "USGS:06928300:00011:00015",
  "USGS:06928300:00011:00001",
  "USGS:06928320:00011:00002",
  "USGS:06928320:00011:00001",
  "USGS:06928330:00011:00004",
  "USGS:06928330:00011:00002",
  "USGS:06928330:00011:00001",
  "USGS:06928359:00011:00002",
  "USGS:06928359:00011:00001",
  "USGS:06928420:00011:00012",
  "USGS:06928420:00011:00002",
  "USGS:06928420:00011:00013",
  "USGS:06929900:00011:00002",
  "USGS:06929900:00011:00001",
  "USGS:06930000:00011:00004",
  "USGS:06930000:00011:00002",
  "USGS:06930000:00011:00014",
  "USGS:06930015:00011:00002",
  "USGS:06930015:00011:00001",
  "USGS:06930060:00011:00013",
  "USGS:06930060:00011:00001",
  "USGS:06932000:00011:00001",
  "USGS:06932000:00011:00007",
  "USGS:06933500:00011:00005",
  "USGS:06933500:00011:00002",
  "USGS:06934000:00011:00004",
  "USGS:06934000:00011:00002",
  "USGS:06934500:00011:00036",
  "USGS:06934500:00011:00003",
  "USGS:06934500:00011:00006",
  "USGS:06934500:00011:00002",
  "USGS:06934500:00011:00037",
  "USGS:06934500:00011:00046",
  "USGS:06934500:00011:00049",
  "USGS:06934500:00011:00039",
  "USGS:06934500:00011:00054",
  "USGS:06934500:00011:00040",
  "USGS:06935450:00011:00012",
  "USGS:06935450:00011:00002",
  "USGS:06935450:00011:00001",
  "USGS:02473000:00011:00020",
  "USGS:02473000:00011:00021",
  "USGS:02473000:00011:00006",
  "USGS:02473000:00011:00005",
  "USGS:02473500:00011:00020",
  "USGS:02473500:00011:00021",
  "USGS:02473500:00011:00004",
  "USGS:02473500:00011:00003",
  "USGS:02474500:00011:00004",
  "USGS:02474500:00011:00003",
  "USGS:02474560:00011:00019",
  "USGS:02474560:00011:00004",
  "USGS:02474560:00011:00003",
  "USGS:02475000:00011:00017",
  "USGS:02475000:00011:00018",
  "USGS:02475000:00011:00004",
  "USGS:02475000:00011:00003",
  "USGS:02475500:00011:00004",
  "USGS:06935850:00011:00005",
  "USGS:06935850:00011:00002",
  "USGS:06935850:00011:00004",
  "USGS:06935890:00011:00015",
  "USGS:06935890:00011:00003",
  "USGS:06935890:00011:00001",
  "USGS:06935955:00011:00002",
  "USGS:06935955:00011:00004",
  "USGS:06935965:00011:00019",
  "USGS:06935965:00011:00020",
  "USGS:06935965:00011:00021",
  "USGS:06935965:00011:00014",
  "USGS:06935965:00011:00002",
  "USGS:06935965:00011:00003",
  "USGS:06935980:00011:00003",
  "USGS:06935980:00011:00002",
  "USGS:06935997:00011:00002",
  "USGS:06935997:00011:00001",
  "USGS:06936475:00011:00015",
  "USGS:06936475:00011:00002",
  "USGS:06936475:00011:00005",
  "USGS:06936530:00011:00002",
  "USGS:06936530:00011:00001",
  "USGS:07001910:00011:00002",
  "USGS:07001910:00011:00001",
  "USGS:07001985:00011:00002",
  "USGS:07001985:00011:00001",
  "USGS:07005000:00011:00015",
  "USGS:07005000:00011:00002",
  "USGS:07005000:00011:00001",
  "USGS:07010000:00011:00005",
  "USGS:07010000:00011:00002",
  "USGS:07010022:00011:00002",
  "USGS:07010022:00011:00004",
  "USGS:07010030:00011:00002",
  "USGS:07010030:00011:00001",
  "USGS:07010035:00011:00002",
  "USGS:07010035:00011:00001",
  "USGS:07010040:00011:00001",
  "USGS:07010055:00011:00002",
  "USGS:07010055:00011:00001",
  "USGS:07010061:00011:00002",
  "USGS:07010061:00011:00001",
  "USGS:07010070:00011:00002",
  "USGS:07010070:00011:00001",
  "USGS:07010075:00011:00013",
  "USGS:07010075:00011:00001",
  "USGS:07010082:00011:00001",
  "USGS:07010082:00011:00013",
  "USGS:07010086:00011:00002",
  "USGS:07010086:00011:00001",
  "USGS:07010088:00011:00001",
  "USGS:07010088:00011:00012",
  "USGS:07010090:00011:00002",
  "USGS:07010090:00011:00001",
  "USGS:07010094:00011:00002",
  "USGS:07010094:00011:00001",
  "USGS:07010097:00011:00004",
  "USGS:07010097:00011:00006",
  "USGS:07010180:00011:00002",
  "USGS:07010180:00011:00001",
  "USGS:07010208:00011:00016",
  "USGS:07010208:00011:00002",
  "USGS:07010208:00011:00005",
  "USGS:07010350:00011:00001",
  "USGS:07010350:00011:00002",
  "USGS:07013000:00011:00003",
  "USGS:07013000:00011:00005",
  "USGS:07013000:00011:00002",
  "USGS:07014000:00011:00014",
  "USGS:07014000:00011:00003",
  "USGS:07014000:00011:00002",
  "USGS:07014000:00011:00001",
  "USGS:07014500:00011:00005",
  "USGS:07014500:00011:00002",
  "USGS:07015720:00011:00001",
  "USGS:07015720:00011:00004",
  "USGS:07016500:00011:00003",
  "USGS:07016500:00011:00005",
  "USGS:07016500:00011:00002",
  "USGS:07017020:00011:00001",
  "USGS:07017200:00011:00001",
  "USGS:07017200:00011:00004",
  "USGS:07018100:00011:00003",
  "USGS:07018100:00011:00005",
  "USGS:07018100:00011:00002",
  "USGS:07018500:00011:00003",
  "USGS:07018500:00011:00001",
  "USGS:07018500:00011:00004",
  "USGS:07018500:00011:00016",
  "USGS:07019000:00011:00003",
  "USGS:07019000:00011:00006",
  "USGS:07019000:00011:00002",
  "USGS:07019072:00011:00002",
  "USGS:07019072:00011:00004",
  "USGS:07019120:00011:00003",
  "USGS:07019120:00011:00002",
  "USGS:07019130:00011:00012",
  "USGS:07019130:00011:00001",
  "USGS:07019150:00011:00002",
  "USGS:07019150:00011:00001",
  "USGS:07019175:00011:00003",
  "USGS:07019175:00011:00002",
  "USGS:07019185:00011:00015",
  "USGS:07019185:00011:00002",
  "USGS:07019185:00011:00004",
  "USGS:07019195:00011:00002",
  "USGS:07019195:00011:00001",
  "USGS:07019220:00011:00002",
  "USGS:07019220:00011:00005",
  "USGS:02487500:00011:00005",
  "USGS:02487500:00011:00004",
  "USGS:02487500:00011:00003",
  "USGS:02487900:00011:00002",
  "USGS:02488500:00011:00006",
  "USGS:02488500:00011:00019",
  "USGS:02489000:00011:00005",
  "USGS:02489000:00011:00004",
  "USGS:02489000:00011:00003",
  "USGS:02490500:00011:00006",
  "USGS:02490500:00011:00005",
  "USGS:05506350:00011:00014",
  "USGS:05506350:00011:00001",
  "USGS:05506800:00011:00004",
  "USGS:05506800:00011:00002",
  "USGS:05507600:00011:00005",
  "USGS:05507600:00011:00002",
  "USGS:05507800:00011:00015",
  "USGS:05507800:00011:00004",
  "USGS:05507800:00011:00002",
  "USGS:05507820:00011:00011",
  "USGS:05507820:00011:00012",
  "USGS:05507820:00011:00001",
  "USGS:05508000:00011:00019",
  "USGS:05508000:00011:00006",
  "USGS:05508000:00011:00002",
  "USGS:05508805:00011:00005",
  "USGS:05508805:00011:00002",
  "USGS:05514500:00011:00016",
  "USGS:05514500:00011:00001",
  "USGS:05514500:00011:00003",
  "USGS:05514840:00011:00015",
  "USGS:05514840:00011:00013",
  "USGS:05514840:00011:00001",
  "USGS:05514860:00011:00013",
  "USGS:05514860:00011:00001",
  "USGS:06023500:00011:00001",
  "USGS:06023500:00011:00002",
  "USGS:06023800:00011:00002",
  "USGS:06023800:00011:00001",
  "USGS:06024020:00011:00002",
  "USGS:06024020:00011:00001",
  "USGS:06024450:00011:00006",
  "USGS:06024450:00011:00002",
  "USGS:06024450:00011:00005",
  "USGS:06024540:00011:00002",
  "USGS:06024540:00011:00001",
  "USGS:06024580:00011:00001",
  "USGS:06024580:00011:00003",
  "USGS:06024580:00011:00004",
  "USGS:06025250:00011:00004",
  "USGS:06025250:00011:00002",
  "USGS:06025250:00011:00001",
  "USGS:06025500:00011:00019",
  "USGS:06025500:00011:00002",
  "USGS:06025500:00011:00007",
  "USGS:06025500:00011:00011",
  "USGS:06026210:00011:00001",
  "USGS:06026210:00011:00003",
  "USGS:06026210:00011:00002",
  "USGS:06026420:00011:00003",
  "USGS:06026420:00011:00002",
  "USGS:06026420:00011:00001",
  "USGS:06813000:00011:00012",
  "USGS:06813000:00011:00002",
  "USGS:06813000:00011:00003",
  "USGS:06817700:00011:00015",
  "USGS:06817700:00011:00004",
  "USGS:06817700:00011:00002",
  "USGS:06818000:00011:00020",
  "USGS:06818000:00011:00006",
  "USGS:06818000:00011:00002",
  "USGS:06818000:00011:00021",
  "USGS:06818000:00011:00031",
  "USGS:06818000:00011:00024",
  "USGS:06819500:00011:00003",
  "USGS:06819500:00011:00001",
  "USGS:06820410:00011:00012",
  "USGS:06820410:00011:00002",
  "USGS:06820410:00011:00001",
  "USGS:06820500:00011:00006",
  "USGS:06820500:00011:00002",
  "USGS:06821080:00011:00013",
  "USGS:06821080:00011:00018",
  "USGS:06821080:00011:00001",
  "USGS:06821140:00011:00016",
  "USGS:06821150:00011:00004",
  "USGS:06821150:00011:00002",
  "USGS:06821190:00011:00006",
  "USGS:06821190:00011:00002",
  "USGS:06893000:00011:00004",
  "USGS:06893000:00011:00002",
  "USGS:06893060:00011:00001",
  "USGS:06893150:00011:00006",
  "USGS:06893150:00011:00002",
  "USGS:06893150:00011:00004",
  "USGS:06893400:00011:00015",
  "USGS:06893400:00011:00013",
  "USGS:06893400:00011:00001",
  "USGS:06893500:00011:00004",
  "USGS:06893500:00011:00002",
  "USGS:06893557:00011:00005",
  "USGS:06893557:00011:00002",
  "USGS:06893557:00011:00003",
  "USGS:06893562:00011:00001",
  "USGS:06893562:00011:00032",
  "USGS:06893562:00011:00002",
  "USGS:06893578:00011:00013",
  "USGS:06893578:00011:00001",
  "USGS:06893590:00011:00003",
  "USGS:06893620:00011:00011",
  "USGS:06893620:00011:00005",
  "USGS:06893620:00011:00004",
  "USGS:06893620:00011:00001",
  "USGS:06893620:00011:00002",
  "USGS:06893620:00011:00007",
  "USGS:06893620:00011:00009",
  "USGS:06893620:00011:00010",
  "USGS:06893620:00011:00006",
  "USGS:06893620:00011:00008",
  "USGS:06026500:00011:00001",
  "USGS:06026500:00011:00002",
  "USGS:06026500:00011:00007",
  "USGS:06027600:00011:00003",
  "USGS:06027600:00011:00002",
  "USGS:06027600:00011:00001",
  "USGS:06033000:00011:00001",
  "USGS:06033000:00011:00003",
  "USGS:06036650:00011:00008",
  "USGS:06036650:00011:00002",
  "USGS:07020850:00011:00003",
  "USGS:07020850:00011:00002",
  "USGS:07020850:00011:00008",
  "USGS:07020850:00011:00009",
  "USGS:07020850:00011:00025",
  "USGS:07020850:00011:00010",
  "USGS:07020850:00011:00026",
  "USGS:07020850:00011:00028",
  "USGS:07021000:00011:00001",
  "USGS:07021000:00011:00003",
  "USGS:07021020:00011:00001",
  "USGS:07034000:00011:00002",
  "USGS:07035000:00011:00005",
  "USGS:07035000:00011:00002",
  "USGS:07035800:00011:00004",
  "USGS:07035800:00011:00002",
  "USGS:07036100:00011:00004",
  "USGS:07036100:00011:00002",
  "USGS:07037300:00011:00002",
  "USGS:07037300:00011:00001",
  "USGS:07037500:00011:00004",
  "USGS:07037500:00011:00002",
  "USGS:07039000:00011:00003",
  "USGS:07039000:00011:00002",
  "USGS:07039500:00011:00004",
  "USGS:07039500:00011:00002",
  "USGS:07043500:00011:00001",
  "USGS:07043500:00011:00007",
  "USGS:07050152:00011:00002",
  "USGS:07050152:00011:00001",
  "USGS:07050690:00011:00003",
  "USGS:07050690:00011:00016",
  "USGS:07050690:00011:00001",
  "USGS:07050700:00011:00017",
  "USGS:07050700:00011:00002",
  "USGS:07050700:00011:00005",
  "USGS:07052000:00011:00016",
  "USGS:07052000:00011:00002",
  "USGS:07052000:00011:00005",
  "USGS:07052100:00011:00020",
  "USGS:07052100:00011:00002",
  "USGS:07052100:00011:00006",
  "USGS:07052120:00011:00002",
  "USGS:07052120:00011:00004",
  "USGS:07052152:00011:00002",
  "USGS:07052152:00011:00004",
  "USGS:07052250:00011:00002",
  "USGS:07052250:00011:00007",
  "USGS:07052345:00011:00016",
  "USGS:07052345:00011:00015",
  "USGS:07052345:00011:00001",
  "USGS:07052500:00011:00003",
  "USGS:07052500:00011:00005",
  "USGS:07052500:00011:00002",
  "USGS:07052820:00011:00002",
  "USGS:07052820:00011:00001",
  "USGS:07053450:00011:00001",
  "USGS:07053450:00011:00014",
  "USGS:07053450:00011:00002",
  "USGS:07053600:00011:00004",
  "USGS:07053600:00011:00002",
  "USGS:07053600:00011:00037",
  "USGS:07053600:00011:00005",
  "USGS:07053810:00011:00003",
  "USGS:07053810:00011:00015",
  "USGS:07053810:00011:00001",
  "USGS:07053820:00011:00002",
  "USGS:07053820:00011:00001",
  "USGS:07054080:00011:00002",
  "USGS:07054080:00011:00001",
  "USGS:07057500:00011:00005",
  "USGS:07057500:00011:00002",
  "USGS:07058000:00011:00001",
  "USGS:07058000:00011:00003",
  "USGS:07061270:00011:00017",
  "USGS:07061270:00011:00014",
  "USGS:07061270:00011:00002",
  "USGS:07061270:00011:00001",
  "USGS:07061270:00011:00018",
  "USGS:07061270:00011:00019",
  "USGS:07061270:00011:00021",
  "USGS:07061270:00011:00020",
  "USGS:07061270:00011:00022",
  "USGS:07061290:00011:00016",
  "USGS:07061290:00011:00018",
  "USGS:07061290:00011:00002",
  "USGS:07061290:00011:00001",
  "USGS:07061290:00011:00014",
  "USGS:07061290:00011:00012",
  "USGS:02475500:00011:00003",
  "USGS:07061290:00011:00013",
  "USGS:07061290:00011:00015",
  "USGS:07061290:00011:00017",
  "USGS:07061500:00011:00005",
  "USGS:07061500:00011:00002",
  "USGS:07061600:00011:00003",
  "USGS:07061600:00011:00002",
  "USGS:07061600:00011:00001",
  "USGS:07061900:00011:00016",
  "USGS:07061900:00011:00015",
  "USGS:07061900:00011:00001",
  "USGS:07062000:00011:00004",
  "USGS:07062000:00011:00015",
  "USGS:07062050:00011:00001",
  "USGS:07062500:00011:00002",
  "USGS:07062500:00011:00004",
  "USGS:07062575:00011:00012",
  "USGS:07062575:00011:00002",
  "USGS:07062575:00011:00013",
  "USGS:07063000:00011:00003",
  "USGS:07063000:00011:00006",
  "USGS:07063000:00011:00002",
  "USGS:07064440:00011:00012",
  "USGS:07064440:00011:00002",
  "USGS:07064440:00011:00001",
  "USGS:07064533:00011:00013",
  "USGS:07064533:00011:00001",
  "USGS:07065200:00011:00016",
  "USGS:07065200:00011:00018",
  "USGS:07065200:00011:00015",
  "USGS:07065200:00011:00001",
  "USGS:07065495:00011:00015",
  "USGS:07065495:00011:00002",
  "USGS:07065495:00011:00003",
  "USGS:07066000:00011:00016",
  "USGS:07066000:00011:00001",
  "USGS:07066000:00011:00004",
  "USGS:07067000:00011:00016",
  "USGS:07067000:00011:00004",
  "USGS:07067000:00011:00002",
  "USGS:07067500:00011:00002",
  "USGS:07067500:00011:00016",
  "USGS:06041000:00011:00005",
  "USGS:06041000:00011:00006",
  "USGS:06041000:00011:00002",
  "USGS:06043500:00011:00001",
  "USGS:06043500:00011:00004",
  "USGS:06048650:00011:00002",
  "USGS:06048650:00011:00001",
  "USGS:06052500:00011:00001",
  "USGS:06052500:00011:00007",
  "USGS:06052500:00011:00002",
  "USGS:06054500:00011:00005",
  "USGS:06054500:00011:00006",
  "USGS:06054500:00011:00002",
  "USGS:06061500:00011:00001",
  "USGS:06061500:00011:00003",
  "USGS:06062500:00011:00001",
  "USGS:06062500:00011:00003",
  "USGS:06063000:00011:00001",
  "USGS:02476500:00011:00004",
  "USGS:02476500:00011:00003",
  "USGS:02476600:00011:00004",
  "USGS:02476600:00011:00003",
  "USGS:02477000:00011:00005",
  "USGS:02477000:00011:00004",
  "USGS:02477500:00011:00003",
  "USGS:02478500:00011:00004",
  "USGS:02478500:00011:00003",
  "USGS:02478500:00011:00017",
  "USGS:02479000:00011:00006",
  "USGS:02479000:00011:00005",
  "USGS:02479000:00011:00021",
  "USGS:02479130:00011:00019",
  "USGS:02479130:00011:00004",
  "USGS:02479130:00011:00003",
  "USGS:02479155:00011:00001",
  "USGS:02479155:00011:00019",
  "USGS:02479155:00011:00007",
  "USGS:02479155:00011:00006",
  "USGS:02479300:00011:00008",
  "USGS:02479300:00011:00007",
  "USGS:02479310:00011:00001",
  "USGS:02479310:00011:00003",
  "USGS:02479310:00011:00002",
  "USGS:02479560:00011:00002",
  "USGS:02479560:00011:00003",
  "USGS:0248018020:00011:00001",
  "USGS:02480212:00011:00002",
  "USGS:02480212:00011:00001",
  "USGS:02480212:00011:00003",
  "USGS:02480212:00011:00015",
  "USGS:02480273:00011:00013",
  "USGS:02480273:00011:00001",
  "USGS:02480273:00011:00002",
  "USGS:02480273:00011:00003",
  "USGS:02480285:00011:00003",
  "USGS:02480285:00011:00001",
  "USGS:02480285:00011:00002",
  "USGS:02480285:00011:00013",
  "USGS:02480287:00011:00002",
  "USGS:02480287:00011:00001",
  "USGS:02480287:00011:00003",
  "USGS:02480287:00011:00006",
  "USGS:02481000:00011:00019",
  "USGS:02481000:00011:00005",
  "USGS:02481000:00011:00004",
  "USGS:02481000:00011:00003",
  "USGS:02481270:00011:00002",
  "USGS:02481270:00011:00001",
  "USGS:02481270:00011:00003",
  "USGS:02481270:00011:00023",
  "USGS:02481299:00011:00001",
  "USGS:02481510:00011:00007",
  "USGS:02481510:00011:00006",
  "USGS:02481510:00011:00005",
  "USGS:02481660:00011:00030",
  "USGS:02481661:00011:00003",
  "USGS:02481661:00011:00001",
  "USGS:0248166310:00011:00003",
  "USGS:0248166310:00011:00001",
  "USGS:0248166590:00011:00003",
  "USGS:0248166590:00011:00001",
  "USGS:02481880:00011:00005",
  "USGS:02481880:00011:00004",
  "USGS:02481880:00011:00003",
  "USGS:02482000:00011:00005",
  "USGS:02482000:00011:00018",
  "USGS:02482000:00011:00017",
  "USGS:02482470:00011:00002",
  "USGS:02482470:00011:00001",
  "USGS:02482550:00011:00004",
  "USGS:02482550:00011:00006",
  "USGS:02482550:00011:00005",
  "USGS:02482550:00011:00018",
  "USGS:02483000:00011:00004",
  "USGS:02483000:00011:00006",
  "USGS:02483000:00011:00005",
  "USGS:02483500:00011:00004",
  "USGS:02483500:00011:00003",
  "USGS:02483500:00011:00002",
  "USGS:02484000:00011:00005",
  "USGS:02484000:00011:00004",
  "USGS:02484000:00011:00003",
  "USGS:02484500:00011:00004",
  "USGS:02484500:00011:00006",
  "USGS:02484500:00011:00005",
  "USGS:02484650:00011:00002",
  "USGS:02484650:00011:00001",
  "USGS:02484760:00011:00002",
  "USGS:02484760:00011:00001",
  "USGS:02485498:00011:00003",
  "USGS:02485600:00011:00001",
  "USGS:02485601:00011:00005",
  "USGS:02485700:00011:00005",
  "USGS:02485700:00011:00004",
  "USGS:02485700:00011:00003",
  "USGS:02485800:00011:00003",
  "USGS:02485820:00011:00001",
  "USGS:02485950:00011:00003",
  "USGS:02486000:00011:00019",
  "USGS:02486000:00011:00005",
  "USGS:02486000:00011:00020",
  "USGS:02486100:00011:00004",
  "USGS:02486100:00011:00003",
  "USGS:02486350:00011:00016",
  "USGS:02486350:00011:00001",
  "USGS:06131200:00011:00001",
  "USGS:06131200:00011:00002",
  "USGS:06132000:00011:00016",
  "USGS:06133500:00011:00001",
  "USGS:06133500:00011:00017",
  "USGS:06133500:00011:00004",
  "USGS:06133500:00011:00002",
  "USGS:06133500:00011:00016",
  "USGS:06133500:00011:00019",
  "USGS:06135000:00011:00004",
  "USGS:06135000:00011:00002",
  "USGS:06139500:00011:00004",
  "USGS:06139500:00011:00002",
  "USGS:02437100:00011:00004",
  "USGS:02437100:00011:00011",
  "USGS:02437100:00011:00005",
  "USGS:02437100:00011:00006",
  "USGS:02437100:00011:00007",
  "USGS:02437100:00011:00008",
  "USGS:02437100:00011:00009",
  "USGS:02437100:00011:00010",
  "USGS:02439400:00011:00004",
  "USGS:02439400:00011:00003",
  "USGS:02441300:00011:00002",
  "USGS:02441390:00011:00002",
  "USGS:02441390:00011:00004",
  "USGS:02441390:00011:00005",
  "USGS:02441390:00011:00006",
  "USGS:02441390:00011:00007",
  "USGS:02441390:00011:00008",
  "USGS:02441390:00011:00009",
  "USGS:02443500:00011:00004",
  "USGS:02443500:00011:00003",
  "USGS:02448000:00011:00004",
  "USGS:02448000:00011:00003",
  "USGS:02472000:00011:00004",
  "USGS:02472000:00011:00003",
  "USGS:02472500:00011:00004",
  "USGS:02472500:00011:00003",
  "USGS:02472850:00011:00002",
  "USGS:02472850:00011:00001",
  "USGS:02472980:00011:00001",
  "USGS:06453600:00011:00004",
  "USGS:06453600:00011:00002",
  "USGS:06453600:00011:00003",
  "USGS:06453620:00011:00002",
  "USGS:390750093233401:00011:00002",
  "USGS:390750093233401:00011:00001",
  "USGS:390945091494001:00011:00001",
  "USGS:390945094234001:00011:00001",
  "USGS:391149092072901:00011:00011",
  "USGS:391149092072901:00011:00001",
  "USGS:391222093185501:00011:00001",
  "USGS:391236094170201:00011:00001",
  "USGS:391622093161001:00011:00014",
  "USGS:391622093161001:00011:00013",
  "USGS:391622093161001:00011:00012",
  "USGS:391622093161001:00011:00002",
  "USGS:391622093161001:00011:00015",
  "USGS:391622093161001:00011:00017",
  "USGS:391622093161001:00011:00018",
  "USGS:391622093161001:00011:00001",
  "USGS:391825091285101:00011:00011",
  "USGS:391825091285101:00011:00001",
  "USGS:392045093302401:00011:00001",
  "USGS:392147090541901:00011:00001",
  "USGS:392228094473101:00011:00011",
  "USGS:392228094473101:00011:00001",
  "USGS:392310094154301:00011:00001",
  "USGS:392321092153901:00011:00001",
  "USGS:392954095013101:00011:00005",
  "USGS:392954095013101:00011:00004",
  "USGS:392954095013101:00011:00003",
  "USGS:392954095013101:00011:00002",
  "USGS:392954095013101:00011:00006",
  "USGS:392954095013101:00011:00008",
  "USGS:392954095013101:00011:00009",
  "USGS:392954095013101:00011:00001",
  "USGS:393218095032601:00011:00001",
  "USGS:393544093075601:00011:00001",
  "USGS:393640092303901:00011:00013",
  "USGS:393640092303901:00011:00012",
  "USGS:393640092303901:00011:00011",
  "USGS:393640092303901:00011:00018",
  "USGS:393640092303901:00011:00014",
  "USGS:393640092303901:00011:00016",
  "USGS:393640092303901:00011:00017",
  "USGS:393640092303901:00011:00001",
  "USCE:393810091145600:00011:00001",
  "USGS:394013093400201:00011:00001",
  "USGS:394156092030201:00011:00001",
  "USGS:394201093181101:00011:00001",
  "USGS:394508093132101:00011:00006",
  "USGS:394508093132101:00011:00004",
  "USGS:394508093132101:00011:00003",
  "USGS:394508093132101:00011:00002",
  "USGS:394508093132101:00011:00007",
  "USGS:394508093132101:00011:00005",
  "USGS:394508093132101:00011:00008",
  "USGS:394508093132101:00011:00018",
  "USGS:394508093132101:00011:00001",
  "USGS:395043091262601:00011:00013",
  "USGS:395043091262601:00011:00002",
  "USGS:395355095051601:00011:00001",
  "USGS:400105093591601:00011:00011",
  "USGS:400105093591601:00011:00001",
  "USGS:400251094485901:00011:00002",
  "USGS:400251094485901:00011:00001",
  "USGS:400458093582001:00011:00001",
  "USGS:401057091494501:00011:00001",
  "USGS:401444093442001:00011:00002",
  "USGS:401920092130301:00011:00001",
  "USGS:402657093470201:00011:00011",
  "USGS:402657093470201:00011:00001",
  "USGS:403055094364701:00011:00002",
  "USGS:403301094492301:00011:00011",
  "USGS:403301094492301:00011:00001",
  "USGS:403452092292901:00011:00012",
  "USGS:403452092292901:00011:00002",
  "USGS:403501091420401:00011:00001",
  "USGS:06289000:00011:00001",
  "USGS:06289000:00011:00004",
  "USGS:06294000:00011:00002",
  "USGS:06294000:00011:00009",
  "USGS:06294500:00011:00005",
  "USGS:06294500:00011:00002",
  "USGS:06295000:00011:00002",
  "USGS:06295000:00011:00007",
  "USGS:06295113:00011:00001",
  "USGS:06295113:00011:00004",
  "USGS:06306300:00011:00002",
  "USGS:382726093121601:00011:00001",
  "USGS:382745091275701:00011:00001",
  "USGS:382748093595101:00011:00001",
  "USGS:382836091502301:00011:00001",
  "USGS:383031090384101:00011:00001",
  "USGS:383226092054001:00011:00001",
  "USGS:383302090420201:00011:00011",
  "USGS:383302090420201:00011:00001",
  "USGS:383550092094201:00011:00002",
  "USGS:383628090411901:00011:00001",
  "USGS:383644091124901:00011:00011",
  "USGS:383644091124901:00011:00001",
  "USGS:383906090511401:00011:00001",
  "USGS:383929092464901:00011:00001",
  "USGS:384147093101901:00011:00001",
  "USGS:384258091243001:00011:00002",
  "USGS:384258091243001:00011:00001",
  "USGS:384258092231401:00011:00005",
  "USGS:384258092231401:00011:00004",
  "USGS:384258092231401:00011:00003",
  "USGS:384258092231401:00011:00002",
  "USGS:384258092231401:00011:00006",
  "USGS:384258092231401:00011:00008",
  "USGS:384258092231401:00011:00009",
  "USGS:384258092231401:00011:00001",
  "USGS:384455093201001:00011:00011",
  "USGS:384455093201001:00011:00001",
  "USGS:384534093431101:00011:00001",
  "USGS:384545093331601:00011:00001",
  "USGS:384713091474301:00011:00001",
  "USGS:384737090372001:00011:00001",
  "USGS:384832093192501:00011:00002",
  "USGS:384846090510301:00011:00002",
  "USGS:384849090092001:00011:00003",
  "USGS:384917091594401:00011:00001",
  "USGS:385156092263202:00011:00001",
  "USGS:385428091265001:00011:00002",
  "USGS:385432091343201:00011:00001",
  "USGS:385718092234201:00011:00001",
  "USGS:385837090594701:00011:00001",
  "USGS:385845090583801:00011:00002",
  "USGS:385853092592801:00011:00011",
  "USGS:385853092592801:00011:00001",
  "USGS:390150090542801:00011:00001",
  "USGS:390207092570801:00011:00002",
  "USGS:390651092125101:00011:00001",
  "USGS:01052500:00011:00001",
  "USGS:01052500:00011:00003",
  "USGS:01053500:00011:00020",
  "USGS:01053500:00011:00008",
  "USGS:01053500:00011:00001",
  "USGS:01053500:00011:00005",
  "USGS:01053600:00011:00002",
  "USGS:01053600:00011:00001",
  "USGS:01054000:00011:00001",
  "USGS:01054000:00011:00003",
  "USGS:01054114:00011:00002",
  "USGS:01054114:00011:00001",
  "USGS:010642505:00011:00004",
  "USGS:010642505:00011:00003",
  "USGS:371801093260401:00011:00001",
  "USGS:372022092542201:00011:00001",
  "USGS:372153091322301:00011:00002",
  "USGS:372202094370201:00011:00011",
  "USGS:372202094370201:00011:00001",
  "USGS:372202094370202:00011:00001",
  "USGS:372338094052801:00011:00001",
  "USGS:372521089362401:00011:00011",
  "USGS:372521089362401:00011:00001",
  "USGS:372715090510701:00011:00001",
  "USGS:372853091061801:00011:00001",
  "USGS:372958094161001:00011:00012",
  "USGS:372958094161001:00011:00002",
  "USGS:373056091063801:00011:00001",
  "USGS:373210090180601:00011:00002",
  "USGS:373559090082901:00011:00002",
  "USGS:373620093470301:00011:00001",
  "USGS:373653091330101:00011:00001",
  "USGS:373701093151601:00011:00002",
  "USGS:373905091071001:00011:00001",
  "USGS:373906092385201:00011:00020",
  "USGS:373906092385201:00011:00001",
  "USGS:373955091065901:00011:00012",
  "USGS:373955091065901:00011:00001",
  "USGS:374254094524501:00011:00002",
  "USGS:374649090242601:00011:00001",
  "USGS:375259093181401:00011:00001",
  "USGS:375306090125301:00011:00011",
  "USGS:375306090125301:00011:00001",
  "USCE:375410089511000:00011:00001",
  "USGS:375429092300701:00011:00001",
  "USGS:375617090465401:00011:00002",
  "USGS:375625091480401:00011:00021",
  "USGS:375625091480401:00011:00002",
  "USGS:375749091475001:00011:00002",
  "USGS:375907091432201:00011:00002",
  "USGS:392336094550403:00011:00001",
  "USGS:01073000:00011:00001",
  "USGS:01073000:00011:00003",
  "USGS:01073319:00011:00004",
  "USGS:01073319:00011:00003",
  "USGS:01073319:00011:00002",
  "USGS:01073319:00011:00001",
  "USGS:01073500:00011:00001",
  "USGS:01073500:00011:00003",
  "USGS:010735562:00011:00002",
  "USGS:010735562:00011:00001",
  "USGS:06461500:00011:00020",
  "USGS:06461500:00011:00008",
  "USGS:06461500:00011:00006",
  "USGS:06461500:00011:00007",
  "USGS:06461500:00011:00022",
  "USGS:06461500:00011:00023",
  "USGS:06461500:00011:00024",
  "USGS:06463500:00011:00008",
  "USGS:06463500:00011:00007",
  "USGS:06463720:00011:00001",
  "USGS:06463720:00011:00002",
  "USGS:06465500:00011:00001",
  "USGS:12331500:00011:00021",
  "USGS:07186900:00011:00003",
  "USGS:07186900:00011:00002",
  "USGS:07186900:00011:00001",
  "USGS:07187000:00011:00005",
  "USGS:07187000:00011:00002",
  "USGS:07188653:00011:00012",
  "USGS:07188653:00011:00016",
  "USGS:07188653:00011:00001",
  "USGS:07188838:00011:00001",
  "USGS:07188838:00011:00003",
  "USGS:07188838:00011:00002",
  "USGS:07188885:00011:00003",
  "USGS:07188885:00011:00016",
  "USGS:07188885:00011:00001",
  "USGS:07189000:00011:00015",
  "USGS:07189000:00011:00005",
  "USGS:07189000:00011:00004",
  "USGS:07189100:00011:00015",
  "USGS:07189100:00011:00001",
  "USGS:360252090173201:00011:00001",
  "USGS:360252090173202:00011:00001",
  "USGS:360425089485001:00011:00012",
  "USGS:360425089485001:00011:00002",
  "USGS:361145089394101:00011:00001",
  "USGS:362718089552301:00011:00001",
  "USGS:362955089581801:00011:00002",
  "USGS:363236094290301:00011:00002",
  "USGS:363436092391001:00011:00001",
  "USGS:363442090364301:00011:00002",
  "USGS:363539091384501:00011:00001",
  "USGS:363551090152801:00011:00011",
  "USGS:363551090152801:00011:00001",
  "USGS:363721094173801:00011:00001",
  "USGS:363728093150401:00011:00012",
  "USGS:363728093150401:00011:00001",
  "USGS:363855093134701:00011:00001",
  "USGS:364006093200301:00011:00001",
  "USGS:364059093520001:00011:00001",
  "USGS:364313094121101:00011:00012",
  "USGS:364324091515001:00011:00011",
  "USGS:364324091515001:00011:00001",
  "USGS:364453093543601:00011:00011",
  "USGS:364453093543601:00011:00001",
  "USGS:364453093543602:00011:00001",
  "USGS:364643089212301:00011:00002",
  "USGS:364818094185301:00011:00001",
  "USGS:364818094185302:00011:00012",
  "USGS:364818094185302:00011:00001",
  "USGS:365319089331001:00011:00012",
  "USGS:365319089331001:00011:00002",
  "USGS:365415093342301:00011:00001",
  "USGS:365451093555501:00011:   NA",
  "USGS:365559092030001:00011:00001",
  "USGS:365602092395101:00011:00002",
  "USGS:365602092395101:00011:00001",
  "USGS:365634093542701:00011:00001",
  "USGS:365644094001301:00011:00001",
  "USGS:365645093431601:00011:00002",
  "USGS:365654091001301:00011:00002",
  "USGS:365949091421401:00011:00001",
  "USGS:370005093122401:00011:00001",
  "USGS:06772775:00011:00002",
  "USGS:06772775:00011:00001",
  "USGS:06772898:00011:00002",
  "USGS:06772898:00011:00001",
  "USGS:06773500:00011:00001",
  "USGS:06773500:00011:00002",
  "USGS:06774000:00011:00006",
  "USGS:06774000:00011:00005",
  "USGS:06775500:00011:00018",
  "USGS:06775500:00011:00008",
  "USGS:06775500:00011:00007",
  "USGS:06775900:00011:00019",
  "USGS:06775900:00011:00006",
  "USGS:06775900:00011:00005",
  "USGS:06781600:00011:00012",
  "USGS:06781600:00011:00002",
  "USGS:06781600:00011:00001",
  "USGS:06785000:00011:00001",
  "USGS:06785000:00011:00002",
  "USGS:06785500:00011:00001",
  "USGS:06785500:00011:00002",
  "USGS:06786000:00011:00007",
  "USGS:06786000:00011:00006",
  "USGS:06790500:00011:00001",
  "USGS:06790500:00011:00002",
  "USGS:06790500:00011:00022",
  "USGS:06792500:00011:00005",
  "USGS:06792500:00011:00004",
  "USGS:06793000:00011:00021",
  "USGS:06037500:00011:00001",
  "USGS:06037500:00011:00002",
  "USGS:06037500:00011:00006",
  "USGS:06037500:00011:00003",
  "USGS:06038500:00011:00006",
  "USGS:06038500:00011:00002",
  "USGS:06038500:00011:00003",
  "USGS:06038500:00011:00004",
  "USGS:06038800:00011:00001",
  "USGS:06038800:00011:00002",
  "USGS:06038800:00011:00006",
  "USGS:06040000:00011:00003",
  "USGS:06040000:00011:00001",
  "USGS:06040000:00011:00002",
  "USGS:06040800:00011:00002",
  "USGS:06040800:00011:00001",
  "USGS:09415250:00011:00001",
  "USGS:09415460:00011:00002",
  "USGS:09415460:00011:00001",
  "USGS:09415510:00011:00001",
  "USGS:09415510:00011:00002",
  "USGS:09415558:00011:00002",
  "USGS:09415558:00011:00001",
  "USGS:09415589:00011:00002",
  "USGS:09415589:00011:00001",
  "USGS:09415590:00011:00001",
  "USGS:09415590:00011:00002",
  "USGS:301141089320300:00011:00008",
  "USGS:301141089320300:00011:00001",
  "USGS:301141089320300:00011:00009",
  "USGS:301141089320300:00011:00027",
  "USGS:301429089145600:00011:00002",
  "USGS:301429089145600:00011:00001",
  "USGS:301429089145600:00011:00014",
  "USGS:301429089145600:00011:00024",
  "USGS:301527088521500:00011:00001",
  "USGS:301527088521500:00011:00004",
  "USGS:301527088521500:00011:00002",
  "USGS:301527088521500:00011:00021",
  "USGS:301527088521500:00011:00023",
  "USGS:301527088521500:00011:00020",
  "USGS:301849088350000:00011:00001",
  "USGS:301849088350000:00011:00004",
  "USGS:301849088350000:00011:00002",
  "USGS:301849088350000:00011:00021",
  "USGS:301912088583300:00011:00002",
  "USGS:301912088583300:00011:00001",
  "USGS:301912088583300:00011:00003",
  "USGS:301912088583300:00011:00023",
  "USGS:301912088583300:00011:00021",
  "USGS:301912088583300:00011:00022",
  "USGS:302318088512600:00011:00001",
  "USGS:302318088512600:00011:00013",
  "USGS:302318088512600:00011:00002",
  "USGS:302318088512600:00011:00017",
  "USGS:3109200904830:00011:00001",
  "USGS:314115088392301:00011:00003",
  "USGS:321759088451400:00011:00005",
  "USGS:321759088451400:00011:00001",
  "USGS:321759088451400:00011:00002",
  "USGS:322722089161050:00011:00001",
  "USGS:322831088474900:00011:00001",
  "USGS:323045090484300:00011:00002",
  "USGS:323045090484300:00011:00003",
  "USGS:323047090484401:00011:00002",
  "USGS:323047090484401:00011:00014",
  "USGS:323331088461300:00011:00001",
  "USGS:325728091002701:00011:00002",
  "USGS:325728091002701:00011:00001",
  "USGS:325817090464201:00011:00002",
  "USGS:325817090464201:00011:00014",
  "USGS:325903089232550:00011:00001",
  "USGS:330152090595601:00011:00002",
  "USGS:330152090595601:00011:00001",
  "USGS:330304090210100:00011:00003",
  "USGS:330304090210100:00011:00004",
  "USGS:330304090210100:00011:00001",
  "USGS:330548091055100:00011:00004",
  "USGS:330548091055100:00011:00001",
  "USGS:332348090505301:00011:00002",
  "USGS:332348090505301:00011:00001",
  "USGS:333136090244900:00011:00001",
  "USGS:333136090244900:00011:00007",
  "USGS:333136090244900:00011:00002",
  "USGS:333145090261901:00011:00002",
  "USGS:333145090261901:00011:00001",
  "USGS:333251090323801:00011:00001",
  "USGS:333420090445900:00011:00002",
  "USGS:333420090445900:00011:00003",
  "USGS:333420090445900:00011:00001",
  "USGS:333601090450000:00011:00002",
  "USGS:333601090450000:00011:00003",
  "USGS:333601090450000:00011:00001",
  "USGS:333830090394600:00011:00012",
  "USGS:333830090394600:00011:00002",
  "USGS:333830090394600:00011:00013",
  "USGS:333830090394600:00011:00003",
  "USGS:333830090394600:00011:00001",
  "USGS:333904090123801:00011:00002",
  "USGS:333904090123801:00011:00001",
  "USGS:334215089442701:00011:00002",
  "USGS:334956090402201:00011:00002",
  "USGS:334956090402201:00011:00001",
  "USGS:335054090230200:00011:00003",
  "USGS:335054090230200:00011:00001",
  "USGS:335054090230200:00011:00004",
  "USGS:335911090553901:00011:00001",
  "USGS:341210090343701:00011:00002",
  "USGS:341210090343701:00011:00014",
  "USGS:341404090385600:00011:00021",
  "USGS:341404090385600:00011:00002",
  "USGS:341404090385600:00011:00022",
  "USGS:341404090385600:00011:00003",
  "USGS:341404090385600:00011:00001",
  "USGS:341550090391300:00011:00002",
  "USGS:341550090391300:00011:00003",
  "USGS:341550090391300:00011:00001",
  "USGS:06805600:00011:00001",
  "USGS:06806500:00011:00005",
  "USGS:06806500:00011:00003",
  "USGS:06807000:00011:00006",
  "USGS:06807000:00011:00024",
  "USGS:06807000:00011:00032",
  "USGS:06807000:00011:00047",
  "USGS:06807000:00011:00049",
  "USGS:06807000:00011:00001",
  "USGS:06807000:00011:00002",
  "USGS:06807000:00011:00025",
  "USGS:06807000:00011:00026",
  "USGS:06807000:00011:00027",
  "USGS:06807000:00011:00028",
  "USGS:06807000:00011:00034",
  "USGS:06810070:00011:00002",
  "USGS:06811500:00011:00018",
  "USGS:06811500:00011:00004",
  "USGS:06811500:00011:00003",
  "USGS:06813500:00011:00003",
  "USGS:06813500:00011:00004",
  "USGS:06813500:00011:00002",
  "USGS:06814500:00011:00001",
  "USGS:06814500:00011:00003",
  "USGS:06815000:00011:00001",
  "USGS:06815000:00011:00002",
  "USGS:06821500:00011:00007",
  "USGS:06821500:00011:00006",
  "USGS:06793000:00011:00018",
  "USGS:06794000:00011:00005",
  "USGS:06794650:00011:00002",
  "USGS:06794650:00011:00001",
  "USGS:06795500:00011:00019",
  "USGS:06795500:00011:00004",
  "USGS:06795500:00011:00003",
  "USGS:06795500:00011:00021",
  "USGS:06795500:00011:00020",
  "USGS:06795500:00011:00022",
  "USGS:06796000:00011:00007",
  "USGS:06796000:00011:00006",
  "USGS:06796500:00011:00002",
  "USGS:06796500:00011:00001",
  "USGS:06796550:00011:00002",
  "USGS:06796550:00011:00015",
  "USGS:06796550:00011:00001",
  "USGS:06797500:00011:00005",
  "USGS:06797500:00011:00004",
  "USGS:06799000:00011:00001",
  "USGS:06799000:00011:00002",
  "USGS:06799080:00011:00002",
  "USGS:06799100:00011:00005",
  "USGS:06799100:00011:00004",
  "USGS:06799315:00011:00002",
  "USGS:06799315:00011:00001",
  "USGS:06799315:00011:00015",
  "USGS:06799350:00011:00020",
  "USGS:06799350:00011:00001",
  "USGS:06799350:00011:00002",
  "USGS:06799445:00011:00013",
  "USGS:06799445:00011:00014",
  "USGS:06799500:00011:00004",
  "USGS:06799500:00011:00003",
  "USGS:06799500:00011:00023",
  "USGS:06800000:00011:00027",
  "USGS:06800000:00011:00004",
  "USGS:06800000:00011:00003",
  "USGS:06800500:00011:00019",
  "USGS:06800500:00011:00001",
  "USGS:06800500:00011:00002",
  "USGS:06800500:00011:00007",
  "USGS:06800500:00011:00008",
  "USGS:06800500:00011:00029",
  "USGS:06801000:00011:00004",
  "USGS:06801000:00011:00003",
  "USGS:06801000:00011:00014",
  "USGS:06803000:00011:00005",
  "USGS:06803000:00011:00004",
  "USGS:06803000:00011:00003",
  "USGS:06803080:00011:00016",
  "USGS:06803080:00011:00014",
  "USGS:06803080:00011:00002",
  "USGS:06803080:00011:00001",
  "USGS:06803093:00011:00014",
  "USGS:06803093:00011:00002",
  "USGS:06803093:00011:00001",
  "USGS:06803170:00011:00014",
  "USGS:06803170:00011:00002",
  "USGS:06803170:00011:00001",
  "USGS:06803300:00011:00003",
  "USGS:06803300:00011:00001",
  "USGS:06803300:00011:00002",
  "USGS:06803486:00011:00003",
  "USGS:06803486:00011:00002",
  "USGS:06803486:00011:00001",
  "USGS:06803495:00011:00001",
  "USGS:06803495:00011:00002",
  "USGS:06803500:00011:00003",
  "USGS:06803500:00011:00001",
  "USGS:06803500:00011:00002",
  "USGS:06803502:00011:00002",
  "USGS:06803510:00011:00005",
  "USGS:06803510:00011:00004",
  "USGS:06803513:00011:00002",
  "USGS:06803513:00011:00001",
  "USGS:06803520:00011:00004",
  "USGS:06803520:00011:00003",
  "USGS:06803530:00011:00007",
  "USGS:06803530:00011:00006",
  "USGS:06803555:00011:00001",
  "USGS:06803555:00011:00002",
  "USGS:06804000:00011:00001",
  "USGS:06804000:00011:00002",
  "USGS:06804000:00011:00005",
  "USGS:06804700:00011:00004",
  "USGS:06804700:00011:00003",
  "USGS:06805000:00011:00008",
  "USGS:06805000:00011:00002",
  "USGS:06805000:00011:00003",
  "USGS:06805000:00011:00004",
  "USGS:06805000:00011:00007",
  "USGS:06805020:00011:00001",
  "USGS:06805500:00011:00022",
  "USGS:06805500:00011:00001",
  "USGS:06805500:00011:00002",
  "USGS:06805500:00011:00004",
  "USGS:06805500:00011:00023",
  "USGS:06805500:00011:00024",
  "USGS:06805500:00011:00011",
  "USGS:06805500:00011:00026",
  "USGS:06805570:00011:00001",
  "USGS:405315098304302:00011:00001",
  "USGS:405435098432601:00011:00004",
  "USGS:405435098432601:00011:00003",
  "USGS:405435098432601:00011:00005",
  "USGS:405435098432601:00011:00002",
  "USGS:405435098432601:00011:00009",
  "USGS:405435098432601:00011:00006",
  "USGS:405435098432601:00011:00010",
  "USGS:405435098432601:00011:00011",
  "USGS:405435098432601:00011:00012",
  "USGS:405435098432601:00011:00013",
  "USGS:405435098432601:00011:00014",
  "USGS:405435098432601:00011:00015",
  "USGS:405435098432601:00011:00016",
  "USGS:405435098432601:00011:00017",
  "USGS:405435098432601:00011:00018",
  "USGS:06465500:00011:00008",
  "USGS:06465500:00011:00007",
  "USGS:06465500:00011:00003",
  "USGS:06465500:00011:00023",
  "USGS:06465500:00011:00024",
  "USGS:06465700:00011:00014",
  "USGS:06465700:00011:00002",
  "USGS:06465700:00011:00001",
  "USGS:06466000:00011:00002",
  "USGS:06466000:00011:00013",
  "USGS:06466010:00011:00001",
  "USGS:06466400:00011:00002",
  "USGS:06466400:00011:00001",
  "USGS:06466500:00011:00001",
  "USGS:06466500:00011:00002",
  "USGS:06478523:00011:00001",
  "USGS:06478526:00011:00001",
  "USGS:06486000:00011:00018",
  "USGS:06486000:00011:00001",
  "USGS:06486000:00011:00002",
  "USGS:06600900:00011:00002",
  "USGS:06600900:00011:00001",
  "USGS:06601000:00011:00005",
  "USGS:06601000:00011:00004",
  "USGS:06601200:00011:00002",
  "USGS:06601200:00011:00031",
  "USGS:06601200:00011:00004",
  "USGS:06601200:00011:00003",
  "USGS:06601200:00011:00017",
  "USGS:06601200:00011:00018",
  "USGS:06601200:00011:00019",
  "USGS:06601200:00011:00020",
  "USGS:06609100:00011:00001",
  "USGS:06610000:00011:00024",
  "USGS:06610000:00011:00001",
  "USGS:06610000:00011:00002",
  "USGS:06610705:00011:00003",
  "USGS:06610705:00011:00002",
  "USGS:06610710:00011:00003",
  "USGS:06610710:00011:00002",
  "USGS:06610720:00011:00005",
  "USGS:06610720:00011:00002",
  "USGS:06610720:00011:00001",
  "USGS:06610732:00011:00017",
  "USGS:06610732:00011:00002",
  "USGS:06610732:00011:00001",
  "USGS:06610732:00011:00014",
  "USGS:06610740:00011:00003",
  "USGS:06610740:00011:00002",
  "USGS:06610742:00011:00003",
  "USGS:06610742:00011:00002",
  "USGS:06610750:00011:00020",
  "USGS:06610750:00011:00002",
  "USGS:06610750:00011:00001",
  "USGS:06610750:00011:00016",
  "USGS:06610760:00011:00003",
  "USGS:06610760:00011:00002",
  "USGS:06610765:00011:00005",
  "USGS:06610765:00011:00002",
  "USGS:06610765:00011:00001",
  "USGS:06610770:00011:00020",
  "USGS:06610770:00011:00002",
  "USGS:06610770:00011:00001",
  "USGS:06610773:00011:00003",
  "USGS:06610773:00011:00002",
  "USGS:06610780:00011:00003",
  "USGS:06610780:00011:00002",
  "USGS:06610785:00011:00005",
  "USGS:06610785:00011:00002",
  "USGS:06610785:00011:00001",
  "USGS:06610786:00011:00003",
  "USGS:06610786:00011:00002",
  "USGS:06610788:00011:00003",
  "USGS:06610788:00011:00002",
  "USGS:06610788:00011:00001",
  "USGS:06610793:00011:00005",
  "USGS:06610793:00011:00002",
  "USGS:06610793:00011:00001",
  "USGS:06610795:00011:00003",
  "USGS:06610795:00011:00022",
  "USGS:06610795:00011:00020",
  "USGS:06762500:00011:00001",
  "USGS:06762500:00011:00002",
  "USGS:06764880:00011:00007",
  "USGS:06764880:00011:00006",
  "USGS:06768000:00011:00001",
  "USGS:06768000:00011:00017",
  "USGS:06768000:00011:00002",
  "USGS:06768000:00011:00005",
  "USGS:06768020:00011:00002",
  "USGS:06768020:00011:00001",
  "USGS:06768025:00011:00001",
  "USGS:06768025:00011:00002",
  "USGS:06768035:00011:00002",
  "USGS:06768035:00011:00001",
  "USGS:06769000:00011:00001",
  "USGS:06769000:00011:00002",
  "USGS:06769525:00011:00002",
  "USGS:06769525:00011:00001",
  "USGS:06770200:00011:00001",
  "USGS:06770200:00011:00004",
  "USGS:06770200:00011:00002",
  "USGS:06770200:00011:00005",
  "USGS:06770500:00011:00001",
  "USGS:06770500:00011:00002",
  "USGS:06772100:00011:00014",
  "USGS:06772100:00011:00002",
  "USGS:06772100:00011:00001",
  "USGS:06784000:00011:00001",
  "USGS:06784000:00011:00007",
  "USGS:06784000:00011:00006",
  "USGS:01367690:00011:00002",
  "USGS:01367690:00011:00001",
  "USGS:01367800:00011:00018",
  "USGS:01367800:00011:00007",
  "USGS:01367800:00011:00006",
  "USGS:06306300:00011:00003",
  "USGS:06306300:00011:00004",
  "USGS:06307500:00011:00001",
  "USGS:06307500:00011:00004",
  "USGS:06307500:00011:00002",
  "USGS:06307600:00011:00001",
  "USGS:06307600:00011:00004",
  "USGS:06307600:00011:00003",
  "USGS:06307616:00011:00001",
  "USGS:06307616:00011:00003",
  "USGS:06307616:00011:00005",
  "USGS:06307740:00011:00001",
  "USGS:06307740:00011:00004",
  "USGS:06307740:00011:00002",
  "USGS:06307740:00011:00005",
  "USGS:06307830:00011:00002",
  "USGS:06307830:00011:00010",
  "USGS:06307830:00011:00012",
  "USGS:06308400:00011:00001",
  "USGS:06308400:00011:00004",
  "USGS:06308500:00011:00006",
  "USGS:06308500:00011:00002",
  "USGS:06308500:00011:00008",
  "USGS:06309000:00011:00006",
  "USGS:06309000:00011:00002",
  "USGS:06324500:00011:00002",
  "USGS:06324500:00011:00006",
  "USGS:06324500:00011:00018",
  "USGS:06326500:00011:00006",
  "USGS:06326500:00011:00001",
  "USGS:06327500:00011:00001",
  "USGS:06327500:00011:00006",
  "USGS:06329500:00011:00005",
  "USGS:06329500:00011:00002",
  "USGS:12301300:00011:00002",
  "USGS:12301300:00011:00004",
  "USGS:12301933:00011:00009",
  "USGS:12301933:00011:00008",
  "USGS:12302055:00011:00002",
  "USGS:12302055:00011:00007",
  "USGS:12304500:00011:00002",
  "USGS:12304500:00011:00003",
  "USGS:12323240:00011:00002",
  "USGS:12323240:00011:00003",
  "USGS:12323250:00011:00001",
  "USGS:12323250:00011:00004",
  "USGS:12323600:00011:00002",
  "USGS:12323600:00011:00001",
  "USGS:12323670:00011:00002",
  "USGS:12323670:00011:00001",
  "USGS:12323700:00011:00001",
  "USGS:12323700:00011:00002",
  "USGS:12323700:00011:00004",
  "USGS:12323710:00011:00002",
  "USGS:12323710:00011:00001",
  "USGS:12323720:00011:00002",
  "USGS:12323720:00011:00001",
  "USGS:12323720:00011:00004",
  "USGS:12323750:00011:00003",
  "USGS:12323750:00011:00023",
  "USGS:12323760:00011:00013",
  "USGS:12323760:00011:00002",
  "USGS:12323760:00011:00001",
  "USGS:12323770:00011:00028",
  "USGS:12323770:00011:00001",
  "USGS:12323770:00011:00003",
  "USGS:12323770:00011:00004",
  "USGS:12323800:00011:00002",
  "USGS:12323800:00011:00001",
  "USGS:12323840:00011:00002",
  "USGS:12323840:00011:00001",
  "USGS:12323840:00011:00004",
  "USGS:12323850:00011:00002",
  "USGS:12323850:00011:00001",
  "USGS:12324200:00011:00002",
  "USGS:12324200:00011:00027",
  "USGS:12324400:00011:00002",
  "USGS:12324400:00011:00001",
  "USGS:12324590:00011:00001",
  "USGS:12324590:00011:00020",
  "USGS:12324680:00011:00001",
  "USGS:12324680:00011:00020",
  "USGS:12325000:00011:00001",
  "USGS:12325500:00011:00001",
  "USGS:12325500:00011:00003",
  "USGS:12329500:00011:00001",
  "USGS:12329500:00011:00010",
  "USGS:12330000:00011:00001",
  "USGS:12330000:00011:00003",
  "USGS:12331500:00011:00001",
  "USGS:12331800:00011:00013",
  "USGS:12331800:00011:00001",
  "USGS:12332000:00011:00001",
  "USGS:12332000:00011:00003",
  "USGS:12334510:00011:00023",
  "USGS:12334510:00011:00004",
  "USGS:12334510:00011:00002",
  "USGS:12334550:00011:00001",
  "USGS:12334550:00011:00024",
  "USGS:12335100:00011:00002",
  "USGS:12335100:00011:00001",
  "USGS:12335500:00011:00001",
  "USGS:12335500:00011:00006",
  "USGS:10297010:00011:00001",
  "USGS:10297010:00011:00002",
  "USGS:10297500:00011:00001",
  "USGS:10297500:00011:00002",
  "USGS:10298600:00011:00002",
  "USGS:10298600:00011:00001",
  "USGS:10299100:00011:00001",
  "USGS:10299100:00011:00002",
  "USGS:10300000:00011:00001",
  "USGS:10300000:00011:00002",
  "USGS:10300200:00011:00002",
  "USGS:10300200:00011:00001",
  "USGS:10300600:00011:00001",
  "USGS:10300600:00011:00002",
  "USGS:10301120:00011:00002",
  "USGS:10301120:00011:00001",
  "USGS:10301290:00011:00002",
  "USGS:02490500:00011:00004",
  "USGS:02492110:00011:00003",
  "USGS:02492110:00011:00002",
  "USGS:02492110:00011:00001",
  "USGS:02492343:00011:00002",
  "USGS:02492343:00011:00001",
  "USGS:02492360:00011:00004",
  "USGS:02492360:00011:00003",
  "USGS:02492620:00011:00002",
  "USGS:02492620:00011:00030",
  "USGS:02492620:00011:00028",
  "USGS:02492620:00011:00029",
  "USGS:02492620:00011:00031",
  "USGS:02492620:00011:00001",
  "USGS:02492620:00011:00004",
  "USGS:02492620:00011:00018",
  "USGS:02492620:00011:00016",
  "USGS:02492620:00011:00008",
  "USGS:02492620:00011:00027",
  "USGS:07029270:00011:00002",
  "USGS:07265455:00011:00003",
  "USGS:07265455:00011:00001",
  "USGS:07268000:00011:00004",
  "USGS:07268000:00011:00003",
  "USGS:07274000:00011:00004",
  "USGS:07274000:00011:00003",
  "USGS:07275900:00011:00002",
  "USGS:07275900:00011:00001",
  "USGS:07281600:00011:00013",
  "USGS:07281600:00011:00002",
  "USGS:07281600:00011:00001",
  "USGS:07281600:00011:00019",
  "USGS:07281600:00011:00015",
  "USGS:07282000:00011:00006",
  "USGS:07282000:00011:00003",
  "USGS:07282100:00011:00006",
  "USGS:07283000:00011:00004",
  "USGS:07283000:00011:00003",
  "USGS:07285500:00011:00004",
  "USGS:07285500:00011:00001",
  "USGS:07285500:00011:00014",
  "USGS:07288000:00011:00016",
  "USGS:07288048:00011:00010",
  "USGS:07288048:00011:00011",
  "USGS:07288048:00011:00007",
  "USGS:07288068:00011:00001",
  "USGS:07288280:00011:00002",
  "USGS:07288280:00011:00001",
  "USGS:07288280:00011:00023",
  "USGS:07288500:00011:00003",
  "USGS:07288500:00011:00002",
  "USGS:07288521:00011:00001",
  "USGS:07288580:00011:00005",
  "USGS:07288650:00011:00013",
  "USGS:07288650:00011:00012",
  "USGS:07288650:00011:00001",
  "USGS:07288650:00011:00014",
  "USGS:07288650:00011:00022",
  "USGS:07288650:00011:00031",
  "USGS:07288650:00011:00016",
  "USGS:07288650:00011:00025",
  "USGS:07288700:00011:00013",
  "USGS:07288700:00011:00022",
  "USGS:0728875070:00011:00003",
  "USGS:0728875070:00011:00001",
  "USGS:0728875070:00011:00004",
  "USGS:0728875070:00011:00006",
  "USGS:07288800:00011:00008",
  "USGS:07288800:00011:00003",
  "USGS:07288800:00011:00006",
  "USGS:07288847:00011:00005",
  "USGS:07288847:00011:00003",
  "USGS:07288847:00011:00004",
  "USGS:07288847:00011:00001",
  "USGS:07288847:00011:00017",
  "USGS:07288847:00011:00006",
  "USGS:07288860:00011:00005",
  "USGS:07288860:00011:00003",
  "USGS:07288860:00011:00004",
  "USGS:07288860:00011:00001",
  "USGS:07288860:00011:00017",
  "USGS:07288860:00011:00006",
  "USGS:0728886910:00011:00003",
  "USGS:0728886910:00011:00001",
  "USGS:0728886910:00011:00005",
  "USGS:07288938:00011:00001",
  "USGS:07288939:00011:00007",
  "USGS:07288939:00011:00004",
  "USGS:07288939:00011:00001",
  "USGS:07288955:00011:00005",
  "USGS:07289000:00011:00007",
  "USGS:07289000:00011:00006",
  "USGS:07289000:00011:00005",
  "USGS:07289000:00011:00026",
  "USGS:07289350:00011:00004",
  "USGS:07289350:00011:00003",
  "USGS:07289730:00011:00013",
  "USGS:07290000:00011:00009",
  "USGS:07290000:00011:00008",
  "USGS:07290000:00011:00007",
  "USGS:07290650:00011:00019",
  "USGS:07290650:00011:00018",
  "USGS:07290880:00011:00002",
  "USGS:07291000:00011:00005",
  "USGS:07291000:00011:00008",
  "USGS:07291000:00011:00007",
  "USGS:07292500:00011:00008",
  "USGS:07292500:00011:00007",
  "USGS:07294550:00011:00002",
  "USGS:07294550:00011:00001",
  "USGS:07295000:00011:00005",
  "USGS:07295000:00011:00004",
  "USGS:07295000:00011:00003",
  "USGS:07375280:00011:00002",
  "USGS:07375280:00011:00001",
  "USGS:07376645:00011:00001",
  "USGS:07377385:00011:00001",
  "USGS:301104089253400:00011:00002",
  "USGS:301104089253400:00011:00001",
  "USGS:301104089253400:00011:00003",
  "USGS:301104089253400:00011:00024",
  "USGS:06140500:00011:00002",
  "USGS:06140500:00011:00005",
  "USGS:06142400:00011:00004",
  "USGS:06142400:00011:00002",
  "USGS:06151500:00011:00004",
  "USGS:06151500:00011:00002",
  "USGS:06154100:00011:00005",
  "USGS:06154100:00011:00017",
  "USGS:06154400:00011:00001",
  "USGS:06154400:00011:00003",
  "USGS:06155030:00011:00001",
  "USGS:06155030:00011:00003",
  "USGS:06155500:00011:00001",
  "USGS:06155500:00011:00003",
  "USGS:06164510:00011:00006",
  "USGS:06164510:00011:00002",
  "USGS:06166000:00011:00001",
  "USGS:06167500:00011:00001",
  "USGS:06167500:00011:00002",
  "USGS:06169500:00011:00001",
  "USGS:06169500:00011:00017",
  "USGS:06172310:00011:00002",
  "USGS:06172310:00011:00007",
  "USGS:06174500:00011:00006",
  "USGS:06174500:00011:00002",
  "USGS:06175100:00011:00002",
  "USGS:06175510:00011:00002",
  "USGS:06175520:00011:00001",
  "USGS:06177000:00011:00006",
  "USGS:06177000:00011:00018",
  "USGS:06177500:00011:00001",
  "USGS:06177500:00011:00005",
  "USGS:06177825:00011:00001",
  "USGS:06177825:00011:00003",
  "USGS:06178000:00011:00001",
  "USGS:06178000:00011:00004",
  "USGS:06181000:00011:00001",
  "USGS:06181000:00011:00003",
  "USGS:06183450:00011:00014",
  "USGS:06183450:00011:00001",
  "USGS:06183450:00011:00003",
  "USGS:06185110:00011:00001",
  "USGS:06185110:00011:00002",
  "USGS:06185500:00011:00006",
  "USGS:06185500:00011:00002",
  "USGS:06187915:00011:00002",
  "USGS:06187915:00011:00008",
  "USGS:06187915:00011:00013",
  "USGS:06191000:00011:00002",
  "USGS:06191000:00011:00005",
  "USGS:06191500:00011:00004",
  "USGS:06191500:00011:00002",
  "USGS:06192500:00011:00017",
  "USGS:06192500:00011:00002",
  "USGS:06192500:00011:00007",
  "USGS:06192500:00011:00024",
  "USGS:06192500:00011:00025",
  "USGS:06192500:00011:00026",
  "USGS:06195600:00011:00001",
  "USGS:06195600:00011:00005",
  "USGS:06195750:00011:00001",
  "USGS:06195950:00011:00001",
  "USGS:06200000:00011:00001",
  "USGS:06200000:00011:00003",
  "USGS:06204050:00011:00001",
  "USGS:06204050:00011:00003",
  "USGS:06204070:00011:00004",
  "USGS:06204070:00011:00002",
  "USGS:06204070:00011:00001",
  "USGS:06205000:00011:00013",
  "USGS:06205000:00011:00001",
  "USGS:06205000:00011:00003",
  "USGS:06207500:00011:00002",
  "USGS:06207500:00011:00007",
  "USGS:06208500:00011:00002",
  "USGS:06208500:00011:00007",
  "USGS:06209500:00011:00001",
  "USGS:06209500:00011:00003",
  "USGS:06211000:00011:00001",
  "USGS:06211000:00011:00003",
  "USGS:06211500:00011:00001",
  "USGS:06211500:00011:00003",
  "USGS:06214500:00011:00006",
  "USGS:06214500:00011:00002",
  "USGS:06216900:00011:00001",
  "USGS:06216900:00011:00002",
  "USGS:06287000:00011:00001",
  "USGS:06287000:00011:00002",
  "USGS:06287000:00011:00005",
  "USGS:06287800:00011:00002",
  "USGS:06287800:00011:00001",
  "USGS:06288400:00011:00002",
  "USGS:06288400:00011:00001",
  "USGS:01073587:00011:00004",
  "USGS:01073587:00011:00003",
  "USGS:01073587:00011:00002",
  "USGS:01073587:00011:00001",
  "USGS:01073785:00011:00015",
  "USGS:01073785:00011:00016",
  "USGS:01073785:00011:00002",
  "USGS:01073785:00011:00014",
  "USGS:01074520:00011:00002",
  "USGS:01074520:00011:00003",
  "USGS:01075000:00011:00001",
  "USGS:01075000:00011:00003",
  "USGS:01076000:00011:00001",
  "USGS:01076000:00011:00003",
  "USGS:01076500:00011:00001",
  "USGS:01076500:00011:00003",
  "USGS:01077400:00011:00004",
  "USGS:01077400:00011:00002",
  "USGS:01077400:00011:00001",
  "USGS:01078000:00011:00001",
  "USGS:01078000:00011:00003",
  "USGS:01081000:00011:00001",
  "USGS:01081000:00011:00003",
  "USGS:01081500:00011:00001",
  "USGS:01081500:00011:00003",
  "USGS:01082000:00011:00001",
  "USGS:01082000:00011:00016",
  "USGS:06063000:00011:00002",
  "USGS:06065500:00011:00001",
  "USGS:06065500:00011:00002",
  "USGS:06066500:00011:00015",
  "USGS:06066500:00011:00001",
  "USGS:06066500:00011:00004",
  "USGS:06071300:00011:00002",
  "USGS:06071300:00011:00006",
  "USGS:06073500:00011:00003",
  "USGS:06073500:00011:00001",
  "USGS:06073500:00011:00004",
  "USGS:06074000:00011:00001",
  "USGS:06074000:00011:00002",
  "USGS:06076690:00011:00005",
  "USGS:06076690:00011:00002",
  "USGS:06077200:00011:00003",
  "USGS:06077200:00011:00002",
  "USGS:06077200:00011:00001",
  "USGS:06077500:00011:00003",
  "USGS:06077500:00011:00001",
  "USGS:06077500:00011:00002",
  "USGS:06078200:00011:00005",
  "USGS:06078200:00011:00002",
  "USGS:06078500:00011:00001",
  "USGS:06078500:00011:00003",
  "USGS:06082200:00011:00001",
  "USGS:06082200:00011:00002",
  "USGS:06085800:00011:00005",
  "USGS:06085800:00011:00001",
  "USGS:06085800:00011:00003",
  "USGS:06088500:00011:00002",
  "USGS:06088500:00011:00007",
  "USGS:06089000:00011:00006",
  "USGS:06089000:00011:00002",
  "USGS:06090000:00011:00001",
  "USGS:06090300:00011:00001",
  "USGS:06090300:00011:00004",
  "USGS:06090500:00011:00002",
  "USGS:06090500:00011:00003",
  "USGS:06090650:00011:00002",
  "USGS:06090650:00011:00029",
  "USGS:06090800:00011:00002",
  "USGS:06090800:00011:00007",
  "USGS:06091700:00011:00001",
  "USGS:06091700:00011:00003",
  "USGS:06093200:00011:00001",
  "USGS:06093200:00011:00003",
  "USGS:06099000:00011:00001",
  "USGS:06099000:00011:00003",
  "USGS:06099500:00011:00003",
  "USGS:06099500:00011:00002",
  "USGS:06101500:00011:00002",
  "USGS:06101500:00011:00005",
  "USGS:06102050:00011:00006",
  "USGS:06102050:00011:00001",
  "USGS:06102050:00011:00002",
  "USGS:06102500:00011:00001",
  "USGS:06102500:00011:00004",
  "USGS:06108000:00011:00001",
  "USGS:06108000:00011:00003",
  "USGS:06108800:00011:00002",
  "USGS:06108800:00011:00003",
  "USGS:06109500:00011:00006",
  "USGS:06109500:00011:00002",
  "USGS:06110020:00011:00002",
  "USGS:06110020:00011:00001",
  "USGS:06111800:00011:00003",
  "USGS:06111800:00011:00002",
  "USGS:06114700:00011:00002",
  "USGS:06114700:00011:00001",
  "USGS:06115200:00011:00006",
  "USGS:06115200:00011:00002",
  "USGS:06118500:00011:00001",
  "USGS:06118500:00011:00002",
  "USGS:06119600:00011:00002",
  "USGS:06119600:00011:00001",
  "USGS:06120500:00011:00001",
  "USGS:06120500:00011:00003",
  "USGS:06123030:00011:00002",
  "USGS:06123030:00011:00001",
  "USGS:06125600:00011:00002",
  "USGS:06125600:00011:00001",
  "USGS:06126500:00011:00005",
  "USGS:06126500:00011:00002",
  "USGS:06127500:00011:00001",
  "USGS:06127500:00011:00003",
  "USGS:06130500:00011:00002",
  "USGS:06130500:00011:00003",
  "USGS:06131000:00011:00001",
  "USGS:06131000:00011:00005",
  "USGS:06131000:00011:00002",
  "USGS:01086000:00011:00001",
  "USGS:01086000:00011:00002",
  "USGS:01087000:00011:00005",
  "USGS:01087000:00011:00004",
  "USGS:01087850:00011:00001",
  "USGS:01088400:00011:00003",
  "USGS:01089100:00011:00005",
  "USGS:01089100:00011:00002",
  "USGS:01089100:00011:00003",
  "USGS:01089500:00011:00001",
  "USGS:01089500:00011:00002",
  "USGS:01089925:00011:00002",
  "USGS:01090800:00011:00006",
  "USGS:01090800:00011:00005",
  "USGS:01091000:00011:00004",
  "USGS:01091000:00011:00003",
  "USGS:01091000:00011:00001",
  "USGS:01091000:00011:00002",
  "USGS:01091500:00011:00004",
  "USGS:01091500:00011:00003",
  "USGS:01092000:00011:00001",
  "USGS:01092000:00011:00003",
  "USGS:01093852:00011:00015",
  "USGS:01093852:00011:00014",
  "USGS:01093852:00011:00002",
  "USGS:01093852:00011:00001",
  "USGS:01094000:00011:00001",
  "USGS:01094000:00011:00003",
  "USGS:010642505:00011:00002",
  "USGS:010642505:00011:00001",
  "USGS:01064500:00011:00016",
  "USGS:01064500:00011:00017",
  "USGS:01064500:00011:00004",
  "USGS:01064500:00011:00002",
  "USGS:01064801:00011:00006",
  "USGS:01064801:00011:00002",
  "USGS:01064801:00011:00004",
  "USGS:01072800:00011:00002",
  "USGS:01072800:00011:00001",
  "USGS:01072870:00011:00013",
  "USGS:01072870:00011:00014",
  "USGS:01072870:00011:00002",
  "USGS:01072870:00011:00001",
  "USGS:06454100:00011:00004",
  "USGS:06454100:00011:00002",
  "USGS:06454100:00011:00005",
  "USGS:06454100:00011:00006",
  "USGS:06454100:00011:00007",
  "USGS:12338300:00011:00002",
  "USGS:12338300:00011:00003",
  "USGS:12340000:00011:00035",
  "USGS:12340000:00011:00002",
  "USGS:12340000:00011:00017",
  "USGS:12340500:00011:00002",
  "USGS:12340500:00011:00023",
  "USGS:12342500:00011:00001",
  "USGS:12342500:00011:00003",
  "USGS:12344000:00011:00001",
  "USGS:12344000:00011:00003",
  "USGS:12344000:00011:00002",
  "USGS:12350250:00011:00002",
  "USGS:12350250:00011:00001",
  "USGS:12352500:00011:00015",
  "USGS:12352500:00011:00002",
  "USGS:12352500:00011:00005",
  "USGS:12353000:00011:00002",
  "USGS:12353000:00011:00018",
  "USGS:12354000:00011:00001",
  "USGS:12354000:00011:00005",
  "USGS:12354500:00011:00006",
  "USGS:12354500:00011:00002",
  "USGS:12355500:00011:00025",
  "USGS:12355500:00011:00005",
  "USGS:12355500:00011:00002",
  "USGS:12358500:00011:00004",
  "USGS:12358500:00011:00002",
  "USGS:12359800:00011:00005",
  "USGS:12359800:00011:00002",
  "USGS:12362000:00011:00001",
  "USGS:12362500:00011:00009",
  "USGS:12362500:00011:00008",
  "USGS:12362500:00011:00007",
  "USGS:12363000:00011:00004",
  "USGS:12363000:00011:00005",
  "USGS:12363000:00011:00002",
  "USGS:12363000:00011:00001",
  "USGS:12365700:00011:00002",
  "USGS:12365700:00011:00001",
  "USGS:12366080:00011:00002",
  "USGS:12366080:00011:00001",
  "USGS:12366500:00011:00002",
  "USGS:12366500:00011:00003",
  "USGS:12369000:00011:00005",
  "USGS:12369000:00011:00016",
  "USGS:12369000:00011:00001",
  "USGS:12369000:00011:00017",
  "USGS:12370000:00011:00005",
  "USGS:12370000:00011:00001",
  "USGS:12371550:00011:00002",
  "USGS:12372000:00011:00002",
  "USGS:12372000:00011:00006",
  "USGS:12374250:00011:00001",
  "USGS:12374250:00011:00002",
  "USGS:12375900:00011:00001",
  "USGS:12375900:00011:00005",
  "USGS:12377150:00011:00001",
  "USGS:12377150:00011:00003",
  "USGS:12381400:00011:00001",
  "USGS:12381400:00011:00003",
  "USGS:12388700:00011:00016",
  "USGS:12388700:00011:00001",
  "USGS:12388700:00011:00003",
  "USGS:12389000:00011:00002",
  "USGS:12389000:00011:00005",
  "USGS:12389500:00011:00002",
  "USGS:12389500:00011:00004",
  "USGS:12390700:00011:00001",
  "USGS:12390700:00011:00004",
  "USGS:450524112380701:00011:00001",
  "USGS:453136112420301:00011:00003",
  "USGS:453136112420301:00011:00001",
  "USGS:455024107355601:00011:00001",
  "USGS:462641110561701:00011:00003",
  "USGS:462641110561701:00011:00001",
  "USGS:470709106061401:00011:00001",
  "USGS:472203111112602:00011:00001",
  "USGS:480034105195401:00011:00002",
  "USGS:480608115242901:00011:00002",
  "USGS:480608115242901:00011:00001",
  "USGS:09523800:00011:00001",
  "USGS:09523800:00011:00004",
  "USGS:09525000:00011:00001",
  "USGS:09525000:00011:00002",
  "USGS:09526200:00011:00002",
  "USGS:09526200:00011:00003",
  "USGS:09527590:00011:00013",
  "USGS:09527590:00011:00001",
  "USGS:09527590:00011:00014",
  "USGS:09527594:00011:00003",
  "USGS:09527594:00011:00001",
  "USGS:09527594:00011:00002",
  "USGS:09527597:00011:00003",
  "USGS:09527597:00011:00001",
  "USGS:09527597:00011:00002",
  "USGS:09527630:00011:00003",
  "USGS:09527630:00011:00001",
  "USGS:09527630:00011:00002",
  "USGS:01083000:00011:00008",
  "USGS:01083000:00011:00007",
  "USGS:01085000:00011:00004",
  "USGS:01085000:00011:00003",
  "USGS:01085500:00011:00001",
  "USGS:01085500:00011:00005",
  "USGS:07199450:00011:00002",
  "USGS:07199450:00011:00001",
  "USGS:07202500:00011:00001",
  "USGS:07202500:00011:00002",
  "USGS:07203000:00011:00001",
  "USGS:07203000:00011:00002",
  "USGS:07205500:00011:00002",
  "USGS:07205500:00011:00021",
  "USGS:07206000:00011:00001",
  "USGS:07206000:00011:00002",
  "USGS:07207000:00011:00001",
  "USGS:07207000:00011:00002",
  "USGS:07207500:00011:00001",
  "USGS:07207500:00011:00002",
  "USGS:07208500:00011:00001",
  "USGS:07208500:00011:00002",
  "USGS:07211500:00011:00005",
  "USGS:07211500:00011:00006",
  "USGS:07215500:00011:00001",
  "USGS:07215500:00011:00002",
  "USGS:07216500:00011:00005",
  "USGS:07216500:00011:00006",
  "USGS:07218000:00011:00001",
  "USGS:07218000:00011:00002",
  "USGS:07221500:00011:00005",
  "USGS:07221500:00011:00007",
  "USGS:07226800:00011:00001",
  "USGS:07226800:00011:00014",
  "USGS:07227000:00011:00001",
  "USGS:07227000:00011:00002",
  "USGS:07227100:00011:00001",
  "USGS:07227100:00011:00002",
  "USGS:08253900:00011:00012",
  "USGS:08253900:00011:00002",
  "USGS:08255500:00011:00001",
  "USGS:08255500:00011:00002",
  "USGS:08263500:00011:00001",
  "USGS:08263500:00011:00002",
  "USGS:08265000:00011:00001",
  "USGS:08265000:00011:00002",
  "USGS:08266820:00011:00001",
  "USGS:08266820:00011:00002",
  "USGS:08267500:00011:00001",
  "USGS:08267500:00011:00002",
  "USGS:08269000:00011:00001",
  "USGS:08269000:00011:00002",
  "USGS:363308114553001:00011:00001",
  "USGS:363503115385701:00011:00001",
  "USGS:364650114432001:00011:00001",
  "USGS:364743114533101:00011:00002",
  "USGS:372639114520901:00011:00001",
  "USGS:374215114453101:00011:00002",
  "USGS:380531114534201:00011:00001",
  "USGS:380758115204601:00011:00001",
  "USGS:385521114503601:00011:00001",
  "USGS:390241118513301:00011:00003",
  "USGS:390241118513301:00011:00002",
  "USGS:393310114475001:00011:00002",
  "USGS:394036116183401:00011:00001",
  "USGS:412910117321001:00011:00004",
  "USGS:10308200:00011:00002",
  "USGS:10308200:00011:00003",
  "USGS:10308783:00011:00002",
  "USGS:10308783:00011:00001",
  "USGS:10308784:00011:00002",
  "USGS:10308784:00011:00001",
  "USGS:10308785:00011:00002",
  "USGS:10308785:00011:00001",
  "USGS:103087853:00011:00001",
  "USGS:103087855:00011:00002",
  "USGS:103087855:00011:00001",
  "USGS:103087865:00011:00002",
  "USGS:103087865:00011:00001",
  "USGS:103087889:00011:00002",
  "USGS:103087889:00011:00001",
  "USGS:10308789:00011:00002",
  "USGS:10308789:00011:00001",
  "USGS:103087891:00011:00002",
  "USGS:103087891:00011:00001",
  "USGS:10308794:00011:00001",
  "USGS:10308794:00011:00002",
  "USGS:10310000:00011:00004",
  "USGS:10310000:00011:00003",
  "USGS:01376950:00011:00001",
  "USGS:09415645:00011:00002",
  "USGS:09415645:00011:00001",
  "USGS:09415900:00011:00001",
  "USGS:09415900:00011:00002",
  "USGS:09415908:00011:00002",
  "USGS:09415908:00011:00001",
  "USGS:09415910:00011:00002",
  "USGS:09415910:00011:00001",
  "USGS:09415920:00011:00001",
  "USGS:09415920:00011:00002",
  "USGS:09415927:00011:00002",
  "USGS:09415927:00011:00001",
  "USGS:09416000:00011:00007",
  "USGS:09416000:00011:00001",
  "USGS:09416000:00011:00002",
  "USGS:09417500:00011:00001",
  "USGS:09417500:00011:00002",
  "USGS:09418500:00011:00001",
  "USGS:09418500:00011:00002",
  "USGS:09419000:00011:00001",
  "USGS:09419000:00011:00002",
  "USGS:09419507:00011:00001",
  "USGS:09419507:00011:00002",
  "USGS:09419625:00011:00001",
  "USGS:09419625:00011:00002",
  "USGS:09419659:00011:00003",
  "USGS:09419659:00011:00002",
  "USGS:09419659:00011:00001",
  "USGS:09419665:00011:00003",
  "USGS:09419665:00011:00002",
  "USGS:09419665:00011:00001",
  "USGS:094196781:00011:00003",
  "USGS:094196781:00011:00002",
  "USGS:094196781:00011:00001",
  "USGS:094196784:00011:00003",
  "USGS:094196784:00011:00002",
  "USGS:094196784:00011:00001",
  "USGS:09419679:00011:00002",
  "USGS:09419679:00011:00004",
  "USGS:09419696:00011:00002",
  "USGS:09419696:00011:00001",
  "USGS:09419700:00011:00002",
  "USGS:09419700:00011:00001",
  "USGS:09419740:00011:00003",
  "USGS:09419740:00011:00002",
  "USGS:09419740:00011:00001",
  "USGS:09419745:00011:00003",
  "USGS:09419745:00011:00002",
  "USGS:09419745:00011:00001",
  "USGS:09419753:00011:00002",
  "USGS:09419753:00011:00003",
  "USGS:09419756:00011:00002",
  "USGS:09419756:00011:00001",
  "USGS:09419800:00011:00002",
  "USGS:09419800:00011:00001",
  "USGS:09421500:00011:00017",
  "USGS:09421500:00011:00018",
  "USGS:09421500:00011:00002",
  "USGS:09423000:00011:00002",
  "USGS:09423000:00011:00005",
  "USGS:10243224:00011:00002",
  "USGS:10243224:00011:00001",
  "USGS:102432241:00011:00002",
  "USGS:102432241:00011:00001",
  "USGS:10243260:00011:00001",
  "USGS:10243260:00011:00002",
  "USGS:10243700:00011:00001",
  "USGS:10243700:00011:00002",
  "USGS:10244950:00011:00002",
  "USGS:10244950:00011:00003",
  "USGS:10245100:00011:00002",
  "USGS:10245100:00011:00001",
  "USGS:10245960:00011:00002",
  "USGS:10245960:00011:00001",
  "USGS:10245970:00011:00002",
  "USGS:10245970:00011:00001",
  "USGS:10246835:00011:00001",
  "USGS:10246835:00011:00002",
  "USGS:10249280:00011:00001",
  "USGS:10249280:00011:00003",
  "USGS:10249300:00011:00002",
  "USGS:10249300:00011:00003",
  "USGS:10249300:00011:00004",
  "USGS:10288500:00011:00002",
  "USGS:10288500:00011:00001",
  "USGS:10293048:00011:00002",
  "USGS:10293048:00011:00001",
  "USGS:10293050:00011:00001",
  "USGS:10293050:00011:00002",
  "USGS:10293500:00011:00001",
  "USGS:10293500:00011:00003",
  "USGS:10295000:00011:00001",
  "USGS:10295000:00011:00002",
  "USGS:10297000:00011:00001",
  "USGS:10297000:00011:00005",
  "USGS:422802097031601:00011:00001",
  "USGS:422849099521503:00011:00001",
  "USGS:423148098300601:00011:00002",
  "USGS:423730098560001:00011:00002",
  "USGS:11042400:00011:00001",
  "USGS:11042400:00011:00002",
  "USGS:11042510:00011:00001",
  "USGS:11042510:00011:00002",
  "USGS:11042631:00011:00001",
  "USGS:11042700:00011:00001",
  "USGS:11042800:00011:00002",
  "USGS:11042800:00011:00001",
  "USGS:11042900:00011:00002",
  "USGS:11042900:00011:00001",
  "USGS:11043000:00011:00002",
  "USGS:11044000:00011:00012",
  "USGS:11044000:00011:00001",
  "USGS:11044000:00011:00002",
  "USGS:11044000:00011:00013",
  "USGS:11044000:00011:00014",
  "USGS:11044000:00011:00015",
  "USGS:11044250:00011:00002",
  "USGS:11044250:00011:00001",
  "USGS:10301290:00011:00001",
  "USGS:10301495:00011:00002",
  "USGS:10301495:00011:00001",
  "USGS:10301500:00011:00004",
  "USGS:10301500:00011:00001",
  "USGS:10301500:00011:00002",
  "USGS:10301500:00011:00007",
  "USGS:10301600:00011:00001",
  "USGS:10301600:00011:00002",
  "USGS:10301700:00011:00002",
  "USGS:10301700:00011:00001",
  "USGS:10301720:00011:00002",
  "USGS:10301720:00011:00001",
  "USGS:10301742:00011:00002",
  "USGS:10301742:00011:00001",
  "USGS:10301745:00011:00002",
  "USGS:10301745:00011:00001",
  "USGS:10301755:00011:00004",
  "USGS:10301755:00011:00003",
  "USGS:10302002:00011:00003",
  "USGS:10302002:00011:00002",
  "USGS:10302002:00011:00001",
  "USGS:10302002:00011:00004",
  "USGS:10302025:00011:00004",
  "USGS:10302025:00011:00003",
  "USGS:10308800:00011:00002",
  "USGS:10308800:00011:00004",
  "USGS:10309000:00011:00002",
  "USGS:10309000:00011:00003",
  "USGS:10310400:00011:00001",
  "USGS:10310400:00011:00002",
  "USGS:10310500:00011:00001",
  "USGS:10310500:00011:00002",
  "USGS:10311000:00011:00001",
  "USGS:10311000:00011:00002",
  "USGS:10311100:00011:00001",
  "USGS:10311100:00011:00002",
  "USGS:10311200:00011:00001",
  "USGS:10311200:00011:00002",
  "USGS:10311300:00011:00001",
  "USGS:10311300:00011:00002",
  "USGS:10311400:00011:00001",
  "USGS:10311400:00011:00002",
  "USGS:10312000:00011:00001",
  "USGS:10312000:00011:00002",
  "USGS:10312100:00011:00001",
  "USGS:10312100:00011:00002",
  "USGS:10312150:00011:00002",
  "USGS:10312150:00011:00003",
  "USGS:10312210:00011:00005",
  "USGS:10312210:00011:00002",
  "USGS:10312210:00011:00001",
  "USGS:10312210:00011:00006",
  "USGS:10312275:00011:00001",
  "USGS:10312275:00011:00002",
  "USGS:10313900:00011:00002",
  "USGS:10313900:00011:00001",
  "USGS:10315500:00011:00001",
  "USGS:10315500:00011:00002",
  "USGS:10316500:00011:00001",
  "USGS:10316500:00011:00002",
  "USGS:10317480:00011:00002",
  "USGS:10317480:00011:00001",
  "USGS:10317500:00011:00001",
  "USGS:10317500:00011:00002",
  "USGS:10318500:00011:00001",
  "USGS:10318500:00011:00002",
  "USGS:10319900:00011:00002",
  "USGS:10319900:00011:00001",
  "USGS:10320000:00011:00004",
  "USGS:10320000:00011:00003",
  "USGS:10321000:00011:00002",
  "USGS:10321000:00011:00003",
  "USGS:10321590:00011:00002",
  "USGS:10321590:00011:00001",
  "USGS:10321940:00011:00002",
  "USGS:10321940:00011:00001",
  "USGS:10321950:00011:00002",
  "USGS:10321950:00011:00001",
  "USGS:10322000:00011:00001",
  "USGS:10322000:00011:00002",
  "USGS:10322150:00011:00002",
  "USGS:10322150:00011:00003",
  "USGS:10322500:00011:00003",
  "USGS:10322500:00011:00006",
  "USGS:10322505:00011:00002",
  "USGS:10322505:00011:00001",
  "USGS:103225055:00011:00002",
  "USGS:103225055:00011:00001",
  "USGS:11070465:00011:00001",
  "USGS:10322510:00011:00002",
  "USGS:10322510:00011:00001",
  "USGS:10322535:00011:00002",
  "USGS:10322535:00011:00001",
  "USGS:10322555:00011:00002",
  "USGS:10322555:00011:00001",
  "USGS:10322800:00011:00002",
  "USGS:10322800:00011:00001",
  "USGS:10323425:00011:00002",
  "USGS:10323425:00011:00001",
  "USGS:10324500:00011:00001",
  "USGS:10324500:00011:00002",
  "USGS:10324700:00011:00002",
  "USGS:10324700:00011:00001",
  "USGS:10325000:00011:00001",
  "USGS:10325000:00011:00002",
  "USGS:10327500:00011:00001",
  "USGS:10327500:00011:00002",
  "USGS:10329000:00011:00001",
  "USGS:10329000:00011:00002",
  "USGS:10329500:00011:00001",
  "USGS:10329500:00011:00002",
  "USGS:10333000:00011:00001",
  "USGS:10333000:00011:00002",
  "USGS:10335000:00011:00002",
  "USGS:10335000:00011:00003",
  "USGS:10336698:00011:00003",
  "USGS:10336698:00011:00010",
  "USGS:10336700:00011:00001",
  "USGS:10336700:00011:00002",
  "USGS:10336710:00011:00001",
  "USGS:10336710:00011:00002",
  "USGS:10336730:00011:00001",
  "USGS:10336730:00011:00002",
  "USGS:10347310:00011:00002",
  "USGS:10347310:00011:00005",
  "USGS:10347460:00011:00001",
  "USGS:10347460:00011:00002",
  "USGS:10347460:00011:00005",
  "USGS:10347600:00011:00001",
  "USGS:10347600:00011:00002",
  "USGS:10348000:00011:00001",
  "USGS:10348000:00011:00002",
  "USGS:10348036:00011:00002",
  "USGS:10348036:00011:00001",
  "USGS:10348200:00011:00001",
  "USGS:10348200:00011:00002",
  "USGS:10348200:00011:00006",
  "USGS:10348200:00011:00005",
  "USGS:10348245:00011:00004",
  "USGS:10348245:00011:00002",
  "USGS:10348245:00011:00001",
  "USGS:10348300:00011:00001",
  "USGS:10348300:00011:00002",
  "USGS:10348460:00011:00001",
  "USGS:10348460:00011:00002",
  "USGS:10349300:00011:00001",
  "USGS:10349300:00011:00002",
  "USGS:10349849:00011:00001",
  "USGS:10349849:00011:00002",
  "USGS:10349980:00011:00001",
  "USGS:10349980:00011:00002",
  "USGS:10350000:00011:00001",
  "USGS:10350000:00011:00005",
  "USGS:10350340:00011:00002",
  "USGS:10350340:00011:00001",
  "USGS:10350500:00011:00001",
  "USGS:10350500:00011:00003",
  "USGS:10350500:00011:00008",
  "USGS:10351300:00011:00010",
  "USGS:10351300:00011:00014",
  "USGS:10351400:00011:00001",
  "USGS:10351400:00011:00005",
  "USGS:10351600:00011:00004",
  "USGS:10351600:00011:00001",
  "USGS:10351600:00011:00002",
  "USGS:10351600:00011:00014",
  "USGS:10351650:00011:00002",
  "USGS:10351650:00011:00005",
  "USGS:10351700:00011:00005",
  "USGS:10351700:00011:00001",
  "USGS:10351700:00011:00003",
  "USGS:10351700:00011:00009",
  "USGS:10351700:00011:00002",
  "USGS:10352500:00011:00002",
  "USGS:10352500:00011:00003",
  "USGS:103530001:00011:00001",
  "USGS:103530001:00011:00002",
  "USGS:13105000:00011:00001",
  "USGS:13105000:00011:00002",
  "USGS:13161500:00011:00001",
  "USGS:13161500:00011:00002",
  "USGS:13162225:00011:00002",
  "USGS:13162225:00011:00001",
  "USGS:13174000:00011:00001",
  "USGS:13174000:00011:00002",
  "USGS:13174500:00011:00001",
  "USGS:13174500:00011:00002",
  "USGS:13175100:00011:00002",
  "USGS:13175100:00011:00001",
  "USGS:355906115492601:00011:00002",
  "USGS:355906115492601:00011:00001",
  "USGS:360310115303201:00011:00001",
  "USGS:360956115432801:00011:00001",
  "USGS:362727116013501:00011:00002",
  "USGS:362727116013501:00011:00001",
  "USGS:362727116013502:00011:00002",
  "USGS:11128300:00011:00001",
  "USGS:11128300:00011:00002",
  "USGS:11128500:00011:00001",
  "USGS:11128500:00011:00002",
  "USGS:11129800:00011:00001",
  "USGS:11129800:00011:00002",
  "USGS:11132500:00011:00002",
  "USGS:11132500:00011:00004",
  "USGS:11133000:00011:00003",
  "USGS:11133000:00011:00002",
  "USGS:11133000:00011:00001",
  "USGS:11133000:00011:00004",
  "USGS:11133000:00011:00007",
  "USGS:06823000:00011:00004",
  "USGS:06823000:00011:00003",
  "USGS:06823500:00011:00019",
  "USGS:06823500:00011:00006",
  "USGS:06823500:00011:00005",
  "USGS:06824000:00011:00001",
  "USGS:06824000:00011:00004",
  "USGS:06824500:00011:00001",
  "USGS:06824500:00011:00002",
  "USGS:06827500:00011:00004",
  "USGS:06827500:00011:00003",
  "USGS:06828500:00011:00001",
  "USGS:06828500:00011:00002",
  "USGS:06828500:00011:00018",
  "USGS:06834000:00011:00001",
  "USGS:06834000:00011:00002",
  "USGS:06835500:00011:00001",
  "USGS:06835500:00011:00003",
  "USGS:06836500:00011:00001",
  "USGS:06836500:00011:00003",
  "USGS:06837000:00011:00006",
  "USGS:06837000:00011:00005",
  "USGS:06838000:00011:00019",
  "USGS:06838000:00011:00002",
  "USGS:06838000:00011:00006",
  "USGS:06843500:00011:00001",
  "USGS:06843500:00011:00002",
  "USGS:06844500:00011:00001",
  "USGS:06844500:00011:00002",
  "USGS:06844500:00011:00005",
  "USGS:06847000:00011:00002",
  "USGS:06847000:00011:00005",
  "USGS:06847500:00011:00007",
  "USGS:06847500:00011:00006",
  "USGS:06849000:00011:00001",
  "USGS:06849000:00011:00002",
  "USGS:06852500:00011:00016",
  "USGS:06852500:00011:00015",
  "USGS:06853020:00011:00001",
  "USGS:06853020:00011:00002",
  "USGS:06880800:00011:00006",
  "USGS:06880800:00011:00005",
  "USGS:06881000:00011:00001",
  "USGS:06881000:00011:00002",
  "USGS:06881380:00011:00016",
  "USGS:06881380:00011:00002",
  "USGS:06881380:00011:00001",
  "USGS:06881380:00011:00015",
  "USGS:06882000:00011:00018",
  "USGS:06882000:00011:00008",
  "USGS:06882000:00011:00007",
  "USGS:06883000:00011:00008",
  "USGS:06883000:00011:00003",
  "USGS:06883000:00011:00007",
  "USGS:06884000:00011:00001",
  "USGS:06884000:00011:00002",
  "USGS:094156395:00011:00002",
  "USGS:094156395:00011:00001",
  "USGS:400155101521302:00011:00002",
  "USGS:10256500:00011:00001",
  "USGS:403235101395501:00011:00002",
  "USGS:403954099152101:00011:00001",
  "USGS:404343099272901:00011:00001",
  "USGS:404513098181201:00011:00001",
  "USGS:404513098181202:00011:00001",
  "USGS:404618098504401:00011:00001",
  "USGS:404706101282201:00011:00002",
  "USGS:404717099460501:00011:00001",
  "USGS:404949099445701:00011:00001",
  "USGS:405014099591001:00011:00001",
  "USGS:405040098384503:00011:00004",
  "USGS:405040098384503:00011:00003",
  "USGS:405040098384503:00011:00005",
  "USGS:405040098384503:00011:00002",
  "USGS:405040098384503:00011:00009",
  "USGS:405040098384503:00011:00010",
  "USGS:405040098384503:00011:00011",
  "USGS:405040098384503:00011:00012",
  "USGS:405040098384503:00011:00013",
  "USGS:405040098384503:00011:00014",
  "USGS:405040098384503:00011:00015",
  "USGS:405040098384503:00011:00016",
  "USGS:405040098384503:00011:00017",
  "USGS:405040098384503:00011:00018",
  "USGS:405040098384503:00011:00019",
  "USGS:405040098384503:00011:00020",
  "USGS:405040098384503:00011:00021",
  "USGS:405040098384503:00011:00022",
  "USGS:405040098384503:00011:00023",
  "USGS:405040098384503:00011:00024",
  "USGS:405040098384503:00011:00025",
  "USGS:405040098384503:00011:00026",
  "USGS:405040098384503:00011:00027",
  "USGS:405040098384503:00011:00028",
  "USGS:405040098384503:00011:00029",
  "USGS:405040098384503:00011:00030",
  "USGS:405040098384503:00011:00001",
  "USGS:405040098384503:00011:00007",
  "USGS:405118099514901:00011:00004",
  "USGS:405118099514901:00011:00003",
  "USGS:405118099514901:00011:00005",
  "USGS:405118099514901:00011:00002",
  "USGS:405118099514901:00011:00009",
  "USGS:405118099514901:00011:00006",
  "USGS:405118099514901:00011:00011",
  "USGS:405118099514901:00011:00012",
  "USGS:405118099514901:00011:00013",
  "USGS:405118099514901:00011:00014",
  "USGS:405118099514901:00011:00016",
  "USGS:405118099514901:00011:00017",
  "USGS:405118099514901:00011:00018",
  "USGS:405118099514901:00011:00019",
  "USGS:405118099514901:00011:00021",
  "USGS:405118099514901:00011:00022",
  "USGS:405118099514901:00011:00023",
  "USGS:405118099514901:00011:00024",
  "USGS:405118099514901:00011:00001",
  "USGS:405118099514901:00011:00007",
  "USGS:405129099090201:00011:00001",
  "USGS:405137099085201:00011:00001",
  "USGS:405227098165601:00011:00001",
  "USGS:07075280:00011:00003",
  "USGS:07075280:00011:00006",
  "USGS:07075280:00011:00001",
  "USGS:11452600:00011:00002",
  "USGS:11452600:00011:00001",
  "USGS:11452600:00011:00008",
  "USGS:11452600:00011:00007",
  "USGS:11452800:00011:00003",
  "USGS:11452800:00011:00002",
  "USGS:11452800:00011:00001",
  "USGS:11452800:00011:00006",
  "USGS:11452900:00011:00006",
  "USGS:11452900:00011:00002",
  "USGS:11452900:00011:00001",
  "USGS:11452900:00011:00008",
  "USGS:11453000:00011:00002",
  "USGS:11453000:00011:00005",
  "USGS:11453500:00011:00002",
  "USGS:11453500:00011:00005",
  "USGS:11454000:00011:00002",
  "USGS:11454000:00011:00003",
  "USGS:11455139:00011:00002",
  "USGS:11455139:00011:00003",
  "USGS:09527630:00011:00008",
  "USGS:09527660:00011:00003",
  "USGS:09527660:00011:00001",
  "USGS:09527660:00011:00002",
  "USGS:09527660:00011:00008",
  "USGS:09527700:00011:00004",
  "USGS:09527700:00011:00003",
  "USGS:09527700:00011:00001",
  "USGS:09527700:00011:00002",
  "USGS:09527700:00011:00005",
  "USGS:09530000:00011:00001",
  "USGS:09530000:00011:00005",
  "USGS:09530500:00011:00001",
  "USGS:09530500:00011:00002",
  "USGS:10251290:00011:00002",
  "USGS:10251290:00011:00001",
  "USGS:10251300:00011:00002",
  "USGS:10251300:00011:00001",
  "USGS:10251330:00011:00002",
  "USGS:10251330:00011:00001",
  "USGS:10251330:00011:00003",
  "USGS:10251335:00011:00002",
  "USGS:10251335:00011:00001",
  "USGS:10254005:00011:00001",
  "USGS:10254050:00011:00001",
  "USGS:10254050:00011:00002",
  "USGS:10254970:00011:00002",
  "USGS:10254970:00011:00004",
  "USGS:10255550:00011:00001",
  "USGS:10255550:00011:00002",
  "USGS:10256500:00011:00002",
  "USGS:10257500:00011:00001",
  "USGS:10257500:00011:00002",
  "USGS:10257548:00011:00001",
  "USGS:10257548:00011:00002",
  "USGS:10257549:00011:00001",
  "USGS:10257549:00011:00002",
  "USGS:10257600:00011:00001",
  "USGS:10257600:00011:00002",
  "USGS:10257720:00011:00002",
  "USGS:10257720:00011:00001",
  "USGS:10258000:00011:00001",
  "USGS:10258000:00011:00002",
  "USGS:10258500:00011:00001",
  "USGS:10258500:00011:00002",
  "USGS:10259000:00011:00001",
  "USGS:10259000:00011:00002",
  "USGS:10259050:00011:00001",
  "USGS:10259100:00011:00002",
  "USGS:10259100:00011:00001",
  "USGS:10259200:00011:00001",
  "USGS:10259200:00011:00002",
  "USGS:10259300:00011:00001",
  "USGS:10259300:00011:00002",
  "USGS:10259540:00011:00002",
  "USGS:10260500:00011:00012",
  "USGS:10260500:00011:00001",
  "USGS:10260500:00011:00002",
  "USGS:10260500:00011:00013",
  "USGS:10260500:00011:00014",
  "USGS:10260855:00011:00002",
  "USGS:10260855:00011:00001",
  "USGS:10260950:00011:00003",
  "USGS:10260950:00011:00002",
  "USGS:10260950:00011:00001",
  "USGS:10260950:00011:00004",
  "USGS:10260950:00011:00005",
  "USGS:10261500:00011:00001",
  "USGS:10261500:00011:00002",
  "USGS:10261500:00011:00003",
  "USGS:10261500:00011:00004",
  "USGS:10261500:00011:00020",
  "USGS:10262500:00011:00001",
  "USGS:10262500:00011:00002",
  "USGS:10262500:00011:00090",
  "USGS:10262500:00011:00091",
  "USGS:10263000:00011:00002",
  "USGS:10263500:00011:00002",
  "USGS:10263500:00011:00003",
  "USGS:10265150:00011:00003",
  "USGS:10265150:00011:00002",
  "USGS:10265150:00011:00001",
  "USGS:10265150:00011:00004",
  "USGS:10289500:00011:00002",
  "USGS:10289500:00011:00001",
  "USGS:10290500:00011:00001",
  "USGS:10290500:00011:00002",
  "USGS:10291500:00011:00001",
  "USGS:10291500:00011:00002",
  "USGS:10292500:00011:00001",
  "USGS:10292500:00011:00003",
  "USGS:10293000:00011:00005",
  "USGS:10293000:00011:00004",
  "USGS:10296000:00011:00004",
  "USGS:10296000:00011:00003",
  "USGS:10296500:00011:00001",
  "USGS:10296500:00011:00002",
  "USGS:10296700:00011:00002",
  "USGS:10296750:00011:00001",
  "USGS:10296750:00011:00002",
  "USGS:11274500:00011:00001",
  "USGS:11274500:00011:00002",
  "USGS:11274538:00011:00003",
  "USGS:11274538:00011:00002",
  "USGS:11274538:00011:00001",
  "USGS:11274538:00011:00004",
  "USGS:11274550:00011:00004",
  "USGS:11274550:00011:00002",
  "USGS:11274550:00011:00001",
  "USGS:11274550:00011:00003",
  "USGS:11274630:00011:00001",
  "USGS:11274630:00011:00002",
  "USGS:11274790:00011:00010",
  "USGS:11274790:00011:00009",
  "USGS:11274790:00011:00008",
  "USGS:11274790:00011:00021",
  "USGS:11274790:00011:00011",
  "USGS:11275500:00011:00001",
  "USGS:11275500:00011:00002",
  "USGS:11276500:00011:00001",
  "USGS:11276500:00011:00002",
  "USGS:010965852:00011:00002",
  "USGS:010965852:00011:00003",
  "USGS:01100505:00011:00003",
  "USGS:01100505:00011:00002",
  "USGS:01100505:00011:00001",
  "USGS:01100561:00011:00003",
  "USGS:01100561:00011:00021",
  "USGS:01100561:00011:00001",
  "USGS:01129200:00011:00004",
  "USGS:01129200:00011:00001",
  "USGS:01129200:00011:00003",
  "USGS:01129500:00011:00004",
  "USGS:01129500:00011:00001",
  "USGS:01129500:00011:00003",
  "USGS:01130000:00011:00004",
  "USGS:01130000:00011:00001",
  "USGS:01130000:00011:00005",
  "USGS:01131500:00011:00001",
  "USGS:01131500:00011:00005",
  "USGS:01137500:00011:00001",
  "USGS:01137500:00011:00003",
  "USGS:01144500:00011:00001",
  "USGS:01144500:00011:00003",
  "USGS:01152500:00011:00001",
  "USGS:01152500:00011:00005",
  "USGS:01154500:00011:00002",
  "USGS:01154500:00011:00005",
  "USGS:01154950:00011:00002",
  "USGS:01154950:00011:00001",
  "USGS:01157000:00011:00001",
  "USGS:01157000:00011:00002",
  "USGS:01158000:00011:00001",
  "USGS:01158000:00011:00007",
  "USGS:01158110:00011:00001",
  "USGS:01158600:00011:00001",
  "USGS:01158600:00011:00007",
  "USGS:01160350:00011:00006",
  "USGS:01160350:00011:00002",
  "USGS:01160350:00011:00005",
  "USGS:01161000:00011:00001",
  "USGS:01161000:00011:00003",
  "USGS:09423350:00011:00001",
  "USGS:09423350:00011:00002",
  "USGS:09427500:00011:00001",
  "USGS:09427500:00011:00003",
  "USGS:09427520:00011:00002",
  "USGS:09427520:00011:00005",
  "USGS:09429000:00011:00001",
  "USGS:09429000:00011:00004",
  "USGS:09429000:00011:00006",
  "USGS:09429000:00011:00018",
  "USGS:09429000:00011:00022",
  "USGS:09429100:00011:00002",
  "USGS:09429100:00011:00006",
  "USGS:09429155:00011:00001",
  "USGS:09429155:00011:00002",
  "USGS:09429180:00011:00001",
  "USGS:09429180:00011:00002",
  "USGS:09429200:00011:00001",
  "USGS:09429200:00011:00002",
  "USGS:09429500:00011:00003",
  "USGS:09429600:00011:00002",
  "USGS:09429600:00011:00005",
  "USGS:09521100:00011:00001",
  "USGS:09521100:00011:00007",
  "USGS:09523000:00011:00001",
  "USGS:09523000:00011:00002",
  "USGS:09523000:00011:00010",
  "USGS:09523200:00011:00001",
  "USGS:09523200:00011:00002",
  "USGS:09523200:00011:00012",
  "USGS:09523400:00011:00001",
  "USGS:09523400:00011:00004",
  "USGS:09523600:00011:00001",
  "USGS:09523600:00011:00004",
  "USGS:430054071382901:00011:00001",
  "USGS:431120071284201:00011:00001",
  "USGS:431540071452801:00011:00001",
  "USGS:444657071074401:00011:00002",
  "USGS:444657071074401:00011:00007",
  "USGS:11337080:00011:00012",
  "USGS:11337080:00011:00005",
  "USGS:11337080:00011:00011",
  "USGS:11337080:00011:00006",
  "USGS:11337190:00011:00019",
  "USGS:11337190:00011:00012",
  "USGS:11337190:00011:00003",
  "USGS:11337190:00011:00011",
  "USGS:11337190:00011:00020",
  "USGS:11337190:00011:00061",
  "USGS:11044300:00011:00002",
  "USGS:11044300:00011:00001",
  "USGS:11044350:00011:00002",
  "USGS:11044350:00011:00001",
  "USGS:11044800:00011:00002",
  "USGS:11044800:00011:00001",
  "USGS:11045300:00011:00002",
  "USGS:11045300:00011:00001",
  "USGS:11045600:00011:00001",
  "USGS:11045600:00011:00002",
  "USGS:11045700:00011:00001",
  "USGS:11045700:00011:00002",
  "USGS:11046000:00011:00002",
  "USGS:11046000:00011:00003",
  "USGS:11046100:00011:00001",
  "USGS:11046100:00011:00002",
  "USGS:11046300:00011:00001",
  "USGS:11046300:00011:00002",
  "USGS:11046360:00011:00002",
  "USGS:11046360:00011:00001",
  "USGS:11046530:00011:00002",
  "USGS:11047300:00011:00002",
  "USGS:11047300:00011:00005",
  "USGS:11048200:00011:00001",
  "USGS:11048200:00011:00002",
  "USGS:11048520:00011:00001",
  "USGS:11048600:00011:00001",
  "USGS:11048600:00011:00002",
  "USGS:11051499:00011:00002",
  "USGS:11051499:00011:00003",
  "USGS:11051502:00011:00001",
  "USGS:11051502:00011:00002",
  "USGS:11055500:00011:00002",
  "USGS:11055500:00011:00003",
  "USGS:11055800:00011:00001",
  "USGS:11055800:00011:00002",
  "USGS:11057500:00011:00001",
  "USGS:11057500:00011:00002",
  "USGS:11058000:00011:00001",
  "USGS:11058000:00011:00002",
  "USGS:11058500:00011:00001",
  "USGS:11058500:00011:00002",
  "USGS:11058600:00011:00001",
  "USGS:11058600:00011:00002",
  "USGS:11059300:00011:00003",
  "USGS:11059300:00011:00004",
  "USGS:11060400:00011:00001",
  "USGS:11060400:00011:00002",
  "USGS:11062000:00011:00001",
  "USGS:11062000:00011:00002",
  "USGS:11062399:00011:00002",
  "USGS:11062399:00011:00001",
  "USGS:11062400:00011:00001",
  "USGS:11062400:00011:00002",
  "USGS:11062450:00011:00001",
  "USGS:11062450:00011:00002",
  "USGS:11062700:00011:00001",
  "USGS:11062700:00011:00002",
  "USGS:11062800:00011:00001",
  "USGS:11062800:00011:00002",
  "USGS:11062820:00011:00001",
  "USGS:11062820:00011:00002",
  "USGS:11063510:00011:00001",
  "USGS:11063510:00011:00002",
  "USGS:11063680:00011:00001",
  "USGS:11063680:00011:00002",
  "USGS:11065000:00011:00001",
  "USGS:11065000:00011:00002",
  "USGS:11066460:00011:00004",
  "USGS:11069500:00011:00001",
  "USGS:11069500:00011:00002",
  "USGS:11070150:00011:00001",
  "USGS:11070210:00011:00002",
  "USGS:11070270:00011:00002",
  "USGS:11070270:00011:00003",
  "USGS:11070365:00011:00001",
  "USGS:11070365:00011:00002",
  "USGS:11164500:00011:00001",
  "USGS:11164500:00011:00002",
  "USGS:11166000:00011:00001",
  "USGS:11166000:00011:00002",
  "USGS:11169025:00011:00001",
  "USGS:11169025:00011:00002",
  "USGS:11169025:00011:00013",
  "USGS:11169500:00011:00001",
  "USGS:11169500:00011:00002",
  "USGS:11169750:00011:00001",
  "USGS:11169750:00011:00002",
  "USGS:11169750:00011:00008",
  "USGS:11169750:00011:00004",
  "USGS:11169750:00011:00007",
  "USGS:11169800:00011:00002",
  "USGS:11169800:00011:00005",
  "USGS:405435098432601:00011:00019",
  "USGS:405435098432601:00011:00020",
  "USGS:405435098432601:00011:00021",
  "USGS:405435098432601:00011:00022",
  "USGS:405435098432601:00011:00023",
  "USGS:405435098432601:00011:00024",
  "USGS:405435098432601:00011:00025",
  "USGS:405435098432601:00011:00026",
  "USGS:405435098432601:00011:00027",
  "USGS:405435098432601:00011:00028",
  "USGS:405435098432601:00011:00029",
  "USGS:405435098432601:00011:00030",
  "USGS:405435098432601:00011:00031",
  "USGS:405435098432601:00011:00032",
  "USGS:405435098432601:00011:00033",
  "USGS:405435098432601:00011:00001",
  "USGS:405435098432601:00011:00007",
  "USGS:405445100074001:00011:00001",
  "USGS:405503098441801:00011:00004",
  "USGS:405503098441801:00011:00003",
  "USGS:405503098441801:00011:00005",
  "USGS:405503098441801:00011:00002",
  "USGS:405503098441801:00011:00009",
  "USGS:405503098441801:00011:00006",
  "USGS:405503098441801:00011:00010",
  "USGS:405503098441801:00011:00011",
  "USGS:405503098441801:00011:00012",
  "USGS:405503098441801:00011:00013",
  "USGS:405503098441801:00011:00014",
  "USGS:405503098441801:00011:00015",
  "USGS:405503098441801:00011:00016",
  "USGS:405503098441801:00011:00017",
  "USGS:405503098441801:00011:00018",
  "USGS:405503098441801:00011:00019",
  "USGS:405503098441801:00011:00020",
  "USGS:405503098441801:00011:00021",
  "USGS:405503098441801:00011:00022",
  "USGS:405503098441801:00011:00023",
  "USGS:405503098441801:00011:00024",
  "USGS:405503098441801:00011:00025",
  "USGS:405503098441801:00011:00026",
  "USGS:405503098441801:00011:00027",
  "USGS:405503098441801:00011:00028",
  "USGS:405503098441801:00011:00029",
  "USGS:405503098441801:00011:00030",
  "USGS:405503098441801:00011:00031",
  "USGS:405503098441801:00011:00032",
  "USGS:405503098441801:00011:00033",
  "USGS:405503098441801:00011:00034",
  "USGS:405503098441801:00011:00035",
  "USGS:405503098441801:00011:00036",
  "USGS:405503098441801:00011:00001",
  "USGS:405503098441801:00011:00007",
  "USGS:405632098373501:00011:00001",
  "USGS:405738099504501:00011:00004",
  "USGS:405738099504501:00011:00003",
  "USGS:405738099504501:00011:00005",
  "USGS:405738099504501:00011:00002",
  "USGS:405738099504501:00011:00009",
  "USGS:405738099504501:00011:00006",
  "USGS:405738099504501:00011:00011",
  "USGS:405738099504501:00011:00012",
  "USGS:405738099504501:00011:00013",
  "USGS:405738099504501:00011:00014",
  "USGS:405738099504501:00011:00015",
  "USGS:405738099504501:00011:00016",
  "USGS:405738099504501:00011:00017",
  "USGS:405738099504501:00011:00018",
  "USGS:405738099504501:00011:00019",
  "USGS:405738099504501:00011:00020",
  "USGS:405738099504501:00011:00021",
  "USGS:405738099504501:00011:00022",
  "USGS:405738099504501:00011:00023",
  "USGS:405738099504501:00011:00024",
  "USGS:405738099504501:00011:00025",
  "USGS:405738099504501:00011:00026",
  "USGS:405738099504501:00011:00027",
  "USGS:405738099504501:00011:00028",
  "USGS:405738099504501:00011:00030",
  "USGS:405738099504501:00011:00031",
  "USGS:405738099504501:00011:00032",
  "USGS:405738099504501:00011:00033",
  "USGS:405738099504501:00011:00034",
  "USGS:405738099504501:00011:00001",
  "USGS:405738099504501:00011:00007",
  "USGS:405855098383001:00011:00004",
  "USGS:405855098383001:00011:00003",
  "USGS:405855098383001:00011:00005",
  "USGS:405855098383001:00011:00002",
  "USGS:405855098383001:00011:00009",
  "USGS:405855098383001:00011:00006",
  "USGS:405855098383001:00011:00010",
  "USGS:405855098383001:00011:00011",
  "USGS:405855098383001:00011:00012",
  "USGS:405855098383001:00011:00013",
  "USGS:405855098383001:00011:00014",
  "USGS:405855098383001:00011:00015",
  "USGS:405855098383001:00011:00016",
  "USGS:405855098383001:00011:00017",
  "USGS:405855098383001:00011:00018",
  "USGS:405855098383001:00011:00019",
  "USGS:405855098383001:00011:00020",
  "USGS:405855098383001:00011:00021",
  "USGS:405855098383001:00011:00022",
  "USGS:405855098383001:00011:00023",
  "USGS:405855098383001:00011:00024",
  "USGS:405855098383001:00011:00025",
  "USGS:405855098383001:00011:00026",
  "USGS:405855098383001:00011:00027",
  "USGS:405855098383001:00011:00028",
  "USGS:405855098383001:00011:00029",
  "USGS:405855098383001:00011:00030",
  "USGS:405855098383001:00011:00031",
  "USGS:405855098383001:00011:00032",
  "USGS:405855098383001:00011:00033",
  "USGS:405855098383001:00011:00001",
  "USGS:405855098383001:00011:00007",
  "USGS:405855100073901:00011:00004",
  "USGS:405855100073901:00011:00003",
  "USGS:405855100073901:00011:00005",
  "USGS:405855100073901:00011:00002",
  "USGS:405855100073901:00011:00009",
  "USGS:405855100073901:00011:00006",
  "USGS:405855100073901:00011:00011",
  "USGS:405855100073901:00011:00012",
  "USGS:405855100073901:00011:00013",
  "USGS:405855100073901:00011:00014",
  "USGS:405855100073901:00011:00015",
  "USGS:405855100073901:00011:00016",
  "USGS:405855100073901:00011:00017",
  "USGS:405855100073901:00011:00018",
  "USGS:405855100073901:00011:00019",
  "USGS:405855100073901:00011:00020",
  "USGS:405855100073901:00011:00021",
  "USGS:405855100073901:00011:00022",
  "USGS:405855100073901:00011:00023",
  "USGS:405855100073901:00011:00024",
  "USGS:405855100073901:00011:00025",
  "USGS:405855100073901:00011:00026",
  "USGS:405855100073901:00011:00027",
  "USGS:405855100073901:00011:00028",
  "USGS:405855100073901:00011:00029",
  "USGS:405855100073901:00011:00030",
  "USGS:405855100073901:00011:00031",
  "USGS:405855100073901:00011:00032",
  "USGS:405855100073901:00011:00033",
  "USGS:405855100073901:00011:00034",
  "USGS:405855100073901:00011:00001",
  "USGS:405855100073901:00011:00007",
  "USGS:410102098374201:00011:00004",
  "USGS:410102098374201:00011:00003",
  "USGS:410102098374201:00011:00005",
  "USGS:410102098374201:00011:00002",
  "USGS:410102098374201:00011:00009",
  "USGS:410102098374201:00011:00006",
  "USGS:410102098374201:00011:00010",
  "USGS:410102098374201:00011:00011",
  "USGS:410102098374201:00011:00012",
  "USGS:410102098374201:00011:00013",
  "USGS:410102098374201:00011:00014",
  "USGS:410102098374201:00011:00015",
  "USGS:410102098374201:00011:00016",
  "USGS:410102098374201:00011:00017",
  "USGS:410102098374201:00011:00018",
  "USGS:410102098374201:00011:00019",
  "USGS:410102098374201:00011:00020",
  "USGS:410102098374201:00011:00022",
  "USGS:410102098374201:00011:00023",
  "USGS:410102098374201:00011:00024",
  "USGS:410102098374201:00011:00025",
  "USGS:410102098374201:00011:00026",
  "USGS:410102098374201:00011:00027",
  "USGS:410102098374201:00011:00028",
  "USGS:410102098374201:00011:00029",
  "USGS:410102098374201:00011:00031",
  "USGS:410102098374201:00011:00032",
  "USGS:410102098374201:00011:00001",
  "USGS:410102098374201:00011:00007",
  "USGS:410154099394701:00011:00001",
  "USGS:410156098442601:00011:00002",
  "USGS:410156098442601:00011:00001",
  "USGS:410333095530101:00011:00001",
  "USGS:410333095530101:00011:00023",
  "USGS:410333095530101:00011:00006",
  "USGS:410333095530101:00011:00002",
  "USGS:410333095530101:00011:00004",
  "USGS:410333095530101:00011:00003",
  "USGS:410333095530101:00011:00005",
  "USGS:410618098113401:00011:00001",
  "USGS:410943097575001:00011:00001",
  "USGS:411005096281502:00011:00001",
  "USGS:411219096010601:00011:00018",
  "USGS:411219096010601:00011:00022",
  "USGS:411219096010601:00011:00019",
  "USGS:411219096010601:00011:00002",
  "USGS:411219096010601:00011:00004",
  "USGS:411219096010601:00011:00006",
  "USGS:411219096010601:00011:00008",
  "USGS:411219096010601:00011:00001",
  "USGS:411219096010601:00011:00003",
  "USGS:411219096010601:00011:00005",
  "USGS:411219096010601:00011:00007",
  "USGS:411219096010601:00011:00021",
  "USGS:411219096010601:00011:00023",
  "USGS:411219096010601:00011:00033",
  "USGS:411219096010601:00011:00034",
  "USGS:411219096010601:00011:00035",
  "USGS:411219096010601:00011:00036",
  "USGS:411219096010601:00011:00037",
  "USGS:411219096010601:00011:00038",
  "USGS:411219096010601:00011:00039",
  "USGS:411219096010601:00011:00040",
  "USGS:411219096010601:00011:00041",
  "USGS:411219096010601:00011:00042",
  "USGS:411219096010601:00011:00048",
  "USGS:411219096010601:00011:00049",
  "USGS:411219096010601:00011:00050",
  "USGS:411219096010601:00011:00051",
  "USGS:411219096010601:00011:00009",
  "USGS:411219096010601:00011:00010",
  "USGS:411219096010601:00011:00017",
  "USGS:411232095584201:00011:00001",
  "USGS:411429095583801:00011:00003",
  "USGS:411429095583801:00011:00006",
  "USGS:411429095583801:00011:00004",
  "USGS:411429095583801:00011:00012",
  "USGS:411429095583801:00011:00011",
  "USGS:411429095583801:00011:00013",
  "USGS:411429095583801:00011:00009",
  "USGS:411429095583801:00011:00001",
  "USGS:411429095583801:00011:00005",
  "USGS:411429095583801:00011:00007",
  "USGS:411429095583801:00011:00008",
  "USGS:411429095583801:00011:00002",
  "USGS:411450095582201:00011:00003",
  "USGS:411450095582201:00011:00006",
  "USGS:411450095582201:00011:00004",
  "USGS:411450095582201:00011:00012",
  "USGS:411450095582201:00011:00011",
  "USGS:411450095582201:00011:00013",
  "USGS:411450095582201:00011:00014",
  "USGS:411450095582201:00011:00009",
  "USGS:411450095582201:00011:00001",
  "USGS:411450095582201:00011:00005",
  "USGS:411450095582201:00011:00007",
  "USGS:411450095582201:00011:00008",
  "USGS:411450095582201:00011:00002",
  "USGS:411504096071601:00011:00001",
  "USGS:411701095570601:00011:00001",
  "USGS:411736096170201:00011:00001",
  "USGS:411738097264301:00011:00002",
  "USGS:411857095545301:00011:00001",
  "USGS:412126095565201:00011:00002",
  "USGS:412126095565201:00011:00003",
  "USGS:412126095565201:00011:00004",
  "USGS:412126095565201:00011:00005",
  "USGS:412126095565201:00011:00006",
  "USGS:412336104022801:00011:00003",
  "USGS:412336104022801:00011:00001",
  "USGS:412522100121201:00011:00002",
  "USGS:412522100121201:00011:00001",
  "USGS:412944103452701:00011:00008",
  "USGS:412944103452701:00011:00005",
  "USGS:413130100531202:00011:00001",
  "USGS:413156098591201:00011:00002",
  "USGS:413216102520201:00011:00002",
  "USGS:413216102520201:00011:00001",
  "USGS:413403096135001:00011:00001",
  "USGS:413455102370701:00011:00003",
  "USGS:413455102370701:00011:00001",
  "USGS:413813103334501:00011:00002",
  "USGS:413813103334501:00011:00001",
  "USGS:413853103532102:00011:00003",
  "USGS:413853103532102:00011:00001",
  "USGS:414107102233801:00011:00008",
  "USGS:414107102233801:00011:00005",
  "USGS:414153103561402:00011:00003",
  "USGS:414153103561402:00011:00001",
  "USGS:414607102263301:00011:00001",
  "USGS:415022096434301:00011:00001",
  "USGS:415118103020903:00011:00003",
  "USGS:415118103020903:00011:00001",
  "USGS:415325103392801:00011:00002",
  "USGS:415325103392801:00011:00001",
  "USGS:415559098005201:00011:00002",
  "USGS:415628103554901:00011:00003",
  "USGS:415628103554901:00011:00001",
  "USGS:415654103420401:00011:00002",
  "USGS:415654103420401:00011:00001",
  "USGS:420006102561201:00011:00002",
  "USGS:420006102561201:00011:00001",
  "USGS:420204101200502:00011:00001",
  "USGS:420301103554802:00011:00003",
  "USGS:420301103554802:00011:00001",
  "USGS:420757104024701:00011:00003",
  "USGS:420757104024701:00011:00001",
  "USGS:421210098402001:00011:00002",
  "USGS:422150097402401:00011:00001",
  "USGS:11466320:00011:00001",
  "USGS:11466320:00011:00002",
  "USGS:11466800:00011:00001",
  "USGS:11466800:00011:00002",
  "USGS:11467000:00011:00001",
  "USGS:11467000:00011:00002",
  "USGS:11467000:00011:00006",
  "USGS:11467000:00011:00003",
  "USGS:11467000:00011:00018",
  "USGS:11467000:00011:00019",
  "USGS:11467000:00011:00023",
  "USGS:11467002:00011:00001",
  "USGS:11467200:00011:00001",
  "USGS:11467200:00011:00002",
  "USGS:11467510:00011:00002",
  "USGS:11467510:00011:00001",
  "USGS:11467553:00011:00001",
  "USGS:11467553:00011:00002",
  "USGS:11467553:00011:00005",
  "USGS:11468000:00011:00002",
  "USGS:11468000:00011:00003",
  "USGS:11468500:00011:00002",
  "USGS:11468500:00011:00003",
  "USGS:11468900:00011:00003",
  "USGS:11468900:00011:00001",
  "USGS:11468900:00011:00002",
  "USGS:103366092:00011:00002",
  "USGS:103366092:00011:00003",
  "USGS:10336610:00011:00001",
  "USGS:10336610:00011:00002",
  "USGS:10336610:00011:00009",
  "USGS:10336610:00011:00021",
  "USGS:10336645:00011:00002",
  "USGS:10336645:00011:00006",
  "USGS:10336660:00011:00002",
  "USGS:10336660:00011:00003",
  "USGS:10336676:00011:00002",
  "USGS:10336676:00011:00009",
  "USGS:10336775:00011:00002",
  "USGS:10336775:00011:00003",
  "USGS:10336780:00011:00001",
  "USGS:10336780:00011:00002",
  "USGS:10336780:00011:00003",
  "USGS:10336780:00011:00021",
  "USGS:10337000:00011:00002",
  "USGS:10337500:00011:00003",
  "USGS:10337500:00011:00015",
  "USGS:10337500:00011:00001",
  "USGS:10337500:00011:00002",
  "USGS:10337500:00011:00014",
  "USGS:10338000:00011:00002",
  "USGS:10338000:00011:00004",
  "USGS:10338400:00011:00002",
  "USGS:10338400:00011:00001",
  "USGS:10338500:00011:00002",
  "USGS:10338500:00011:00001",
  "USGS:10338700:00011:00002",
  "USGS:10338700:00011:00001",
  "USGS:10340300:00011:00001",
  "USGS:10340300:00011:00002",
  "USGS:10340500:00011:00001",
  "USGS:10340500:00011:00002",
  "USGS:10342900:00011:00002",
  "USGS:10342900:00011:00001",
  "USGS:10343000:00011:00002",
  "USGS:10343000:00011:00001",
  "USGS:10343500:00011:00001",
  "USGS:10343500:00011:00002",
  "USGS:10343500:00011:00003",
  "USGS:10343500:00011:00006",
  "USGS:10344300:00011:00001",
  "USGS:10344300:00011:00002",
  "USGS:10344400:00011:00001",
  "USGS:10344400:00011:00002",
  "USGS:10344490:00011:00001",
  "USGS:10344490:00011:00002",
  "USGS:10344500:00011:00002",
  "USGS:10344500:00011:00003",
  "USGS:10344505:00011:00002",
  "USGS:10344505:00011:00001",
  "USGS:10346000:00011:00002",
  "USGS:10346000:00011:00001",
  "USGS:10346000:00011:00016",
  "USGS:11012500:00011:00001",
  "USGS:11012500:00011:00002",
  "USGS:11014000:00011:00001",
  "USGS:11014000:00011:00002",
  "USGS:11015000:00011:00001",
  "USGS:11015000:00011:00002",
  "USGS:11016200:00011:00001",
  "USGS:11016200:00011:00002",
  "USGS:11020600:00011:00001",
  "USGS:11020600:00011:00002",
  "USGS:11022100:00011:00001",
  "USGS:11022100:00011:00002",
  "USGS:11022100:00011:00006",
  "USGS:11022200:00011:00001",
  "USGS:11022200:00011:00002",
  "USGS:11022480:00011:00001",
  "USGS:11022480:00011:00002",
  "USGS:11023000:00011:00001",
  "USGS:11023000:00011:00004",
  "USGS:11023000:00011:00005",
  "USGS:11023000:00011:00007",
  "USGS:11023340:00011:00001",
  "USGS:11023340:00011:00002",
  "USGS:11025500:00011:00001",
  "USGS:11025500:00011:00002",
  "USGS:11027000:00011:00003",
  "USGS:11027000:00011:00001",
  "USGS:11027000:00011:00002",
  "USGS:11028500:00011:00001",
  "USGS:11028500:00011:00002",
  "USGS:11042000:00011:00002",
  "USGS:11042000:00011:00003",
  "USGS:323313117033902:00011:00001",
  "USGS:323313117033903:00011:00001",
  "USGS:323313117033904:00011:00001",
  "USGS:323313117033905:00011:00001",
  "USGS:11070465:00011:00002",
  "USGS:11070500:00011:00001",
  "USGS:11070500:00011:00002",
  "USGS:11071900:00011:00002",
  "USGS:11071900:00011:00001",
  "USGS:11072100:00011:00001",
  "USGS:11072100:00011:00002",
  "USGS:11073300:00011:00001",
  "USGS:11073300:00011:00002",
  "USGS:11073360:00011:00001",
  "USGS:11073360:00011:00002",
  "USGS:11073495:00011:00002",
  "USGS:11074000:00011:00001",
  "USGS:11074000:00011:00002",
  "USGS:11074000:00011:00003",
  "USGS:11074000:00011:00021",
  "USGS:11074000:00011:00023",
  "USGS:11074000:00011:00004",
  "USGS:11075720:00011:00001",
  "USGS:11075800:00011:00002",
  "USGS:11077500:00011:00001",
  "USGS:11077500:00011:00002",
  "USGS:11078000:00011:00002",
  "USGS:11078000:00011:00003",
  "USGS:11085000:00011:00001",
  "USGS:11085000:00011:00002",
  "USGS:11087020:00011:00001",
  "USGS:11087020:00011:00002",
  "USGS:11088500:00011:00001",
  "USGS:11088500:00011:00002",
  "USGS:11089200:00011:00002",
  "USGS:11089200:00011:00001",
  "USGS:11089500:00011:00001",
  "USGS:11089500:00011:00002",
  "USGS:11090400:00011:00002",
  "USGS:11090400:00011:00001",
  "USGS:11090600:00011:00002",
  "USGS:11090600:00011:00001",
  "USGS:11092450:00011:00001",
  "USGS:11092450:00011:00002",
  "USGS:11097000:00011:00001",
  "USGS:11097000:00011:00002",
  "USGS:11098000:00011:00001",
  "USGS:11098000:00011:00002",
  "USGS:11101250:00011:00001",
  "USGS:11101250:00011:00002",
  "USGS:11102300:00011:00001",
  "USGS:11102300:00011:00002",
  "USGS:11106550:00011:00002",
  "USGS:11106550:00011:00007",
  "USGS:11109000:00011:00001",
  "USGS:11109000:00011:00002",
  "USGS:11109550:00011:00001",
  "USGS:11109550:00011:00003",
  "USGS:11109600:00011:00002",
  "USGS:11109600:00011:00003",
  "USGS:11109700:00011:00002",
  "USGS:11109700:00011:00001",
  "USGS:11109800:00011:00003",
  "USGS:11109800:00011:00005",
  "USGS:11111500:00011:00002",
  "USGS:11111500:00011:00003",
  "USGS:11113000:00011:00003",
  "USGS:11113000:00011:00007",
  "USGS:11113500:00011:00003",
  "USGS:11113500:00011:00005",
  "USGS:11114495:00011:00001",
  "USGS:11114495:00011:00002",
  "USGS:11118500:00011:00002",
  "USGS:11118500:00011:00005",
  "USGS:11119500:00011:00001",
  "USGS:11119500:00011:00002",
  "USGS:11119745:00011:00002",
  "USGS:11119745:00011:00005",
  "USGS:11119750:00011:00001",
  "USGS:11119750:00011:00002",
  "USGS:11119940:00011:00001",
  "USGS:11119940:00011:00002",
  "USGS:11120000:00011:00002",
  "USGS:11120000:00011:00005",
  "USGS:11120500:00011:00002",
  "USGS:11120500:00011:00003",
  "USGS:11121900:00011:00001",
  "USGS:11121900:00011:00002",
  "USGS:11122000:00011:00003",
  "USGS:11122000:00011:00002",
  "USGS:11122010:00011:00002",
  "USGS:11122010:00011:00001",
  "USGS:11123000:00011:00001",
  "USGS:11123000:00011:00002",
  "USGS:11123500:00011:00001",
  "USGS:11123500:00011:00002",
  "USGS:11124500:00011:00001",
  "USGS:11124500:00011:00002",
  "USGS:11125600:00011:00012",
  "USGS:11125600:00011:00001",
  "USGS:11125600:00011:00002",
  "USGS:11125600:00011:00013",
  "USGS:11126000:00011:00003",
  "USGS:11126000:00011:00001",
  "USGS:11126000:00011:00002",
  "USGS:11126000:00011:00004",
  "USGS:11126000:00011:00015",
  "USGS:11128250:00011:00001",
  "USGS:11128250:00011:00002",
  "USGS:324318117083103:00011:00001",
  "USGS:324318117083104:00011:00001",
  "USGS:324318117083105:00011:00001",
  "USGS:324416117042001:00011:00001",
  "USGS:324416117042002:00011:00001",
  "USGS:324416117042003:00011:00001",
  "USGS:324416117042004:00011:00001",
  "USGS:324416117042005:00011:00001",
  "USGS:324416117042006:00011:00001",
  "USGS:324641117071501:00011:00001",
  "USGS:324641117071502:00011:00001",
  "USGS:324641117071503:00011:00001",
  "USGS:324641117071504:00011:00001",
  "USGS:324641117071505:00011:00001",
  "USGS:330320117024701:00011:00001",
  "USGS:330320117024702:00011:00001",
  "USGS:330320117024703:00011:00001",
  "USGS:11172175:00011:00001",
  "USGS:11172175:00011:00002",
  "USGS:11172945:00011:00012",
  "USGS:11172945:00011:00002",
  "USGS:11172945:00011:00001",
  "USGS:11172955:00011:00002",
  "USGS:11172955:00011:00001",
  "USGS:11173200:00011:00012",
  "USGS:11173200:00011:00001",
  "USGS:11173200:00011:00002",
  "USGS:11173500:00011:00013",
  "USGS:11173500:00011:00001",
  "USGS:11173500:00011:00002",
  "USGS:11173510:00011:00013",
  "USGS:11173510:00011:00002",
  "USGS:11173510:00011:00001",
  "USGS:11173575:00011:00018",
  "USGS:11173575:00011:00002",
  "USGS:11173575:00011:00001",
  "USGS:11173800:00011:00001",
  "USGS:11173800:00011:00002",
  "USGS:11174000:00011:00018",
  "USGS:11174000:00011:00001",
  "USGS:11174000:00011:00002",
  "USGS:11174600:00011:00001",
  "USGS:11174600:00011:00003",
  "USGS:11176400:00011:00002",
  "USGS:11176400:00011:00005",
  "USGS:11176500:00011:00001",
  "USGS:11176500:00011:00002",
  "USGS:11176500:00011:00005",
  "USGS:11176900:00011:00001",
  "USGS:11176900:00011:00005",
  "USGS:11176900:00011:00002",
  "USGS:11176900:00011:00003",
  "USGS:11176900:00011:00004",
  "USGS:11179000:00011:00001",
  "USGS:11179000:00011:00002",
  "USGS:11179000:00011:00006",
  "USGS:11179100:00011:00001",
  "USGS:11179100:00011:00002",
  "USGS:11180500:00011:00001",
  "USGS:11180500:00011:00002",
  "USGS:11180700:00011:00001",
  "USGS:11180700:00011:00002",
  "USGS:11180825:00011:00002",
  "USGS:11180825:00011:00005",
  "USGS:11180900:00011:00002",
  "USGS:11180900:00011:00001",
  "USGS:11180960:00011:00003",
  "USGS:11180960:00011:00006",
  "USGS:11181000:00011:00001",
  "USGS:11181000:00011:00002",
  "USGS:11181008:00011:00001",
  "USGS:11181008:00011:00002",
  "USGS:11181040:00011:00001",
  "USGS:11181040:00011:00002",
  "USGS:11182500:00011:00001",
  "USGS:11182500:00011:00002",
  "USGS:11185185:00011:00017",
  "USGS:11185185:00011:00007",
  "USGS:11185185:00011:00008",
  "USGS:11185185:00011:00003",
  "USGS:11185185:00011:00004",
  "USGS:11189500:00011:00002",
  "USGS:11189500:00011:00004",
  "USGS:11200800:00011:00001",
  "USGS:11200800:00011:00002",
  "USGS:11203580:00011:00012",
  "USGS:11203580:00011:00001",
  "USGS:11203580:00011:00002",
  "USGS:11203580:00011:00013",
  "USGS:11203580:00011:00014",
  "USGS:11204100:00011:00012",
  "USGS:11204100:00011:00001",
  "USGS:11204100:00011:00002",
  "USGS:11204100:00011:00013",
  "USGS:11204100:00011:00014",
  "USGS:11206820:00011:00003",
  "USGS:11206820:00011:00001",
  "USGS:11206820:00011:00002",
  "USGS:11224000:00011:00002",
  "USGS:11224000:00011:00001",
  "USGS:11224500:00011:00001",
  "USGS:11224500:00011:00002",
  "USGS:11251000:00011:00003",
  "USGS:11251000:00011:00001",
  "USGS:11251000:00011:00002",
  "USGS:11251000:00011:00004",
  "USGS:11253130:00011:00001",
  "USGS:11253130:00011:00002",
  "USGS:11253310:00011:00001",
  "USGS:11253310:00011:00002",
  "USGS:11254000:00011:00003",
  "USGS:11254000:00011:00001",
  "USGS:11254000:00011:00002",
  "USGS:11254000:00011:00004",
  "USGS:11255575:00011:00002",
  "USGS:11255575:00011:00001",
  "USGS:11261100:00011:00006",
  "USGS:11261100:00011:00007",
  "USGS:11261100:00011:00009",
  "USGS:11261100:00011:00008",
  "USGS:11261500:00011:00001",
  "USGS:11261500:00011:00002",
  "USGS:11261500:00011:00004",
  "USGS:11261500:00011:00003",
  "USGS:11262900:00011:00006",
  "USGS:11262900:00011:00007",
  "USGS:11262900:00011:00009",
  "USGS:11262900:00011:00008",
  "USGS:11264500:00011:00004",
  "USGS:11264500:00011:00005",
  "USGS:11264500:00011:00006",
  "USGS:11266500:00011:00001",
  "USGS:11266500:00011:00002",
  "USGS:11273400:00011:00003",
  "USGS:11273400:00011:00002",
  "USGS:11273400:00011:00001",
  "USGS:11273400:00011:00004",
  "USGS:11273400:00011:00005",
  "USGS:11273400:00011:00008",
  "USGS:11273400:00011:00009",
  "USGS:11274000:00011:00006",
  "USGS:11274000:00011:00007",
  "USGS:340130117054905:00011:00001",
  "USGS:340136117033901:00011:00001",
  "USGS:340136117033902:00011:00001",
  "USGS:340136117033903:00011:00001",
  "USGS:340136117033904:00011:00001",
  "USGS:340136117033905:00011:00001",
  "USGS:340248117020901:00011:00001",
  "USGS:340248117020902:00011:00001",
  "USGS:340248117020903:00011:00001",
  "USGS:340248117020904:00011:00001",
  "USGS:340408117165301:00011:00001",
  "USGS:340408117165302:00011:00001",
  "USGS:340408117165303:00011:00001",
  "USGS:340439117173902:00011:00001",
  "USGS:340439117173904:00011:00001",
  "USGS:340439117173905:00011:00001",
  "USGS:340439117173906:00011:00001",
  "USGS:340503117104101:00011:00001",
  "USGS:340503117104102:00011:00001",
  "USGS:340503117104103:00011:00001",
  "USGS:340503117104104:00011:00001",
  "USGS:340503117104105:00011:00001",
  "USGS:340521117212001:00011:00001",
  "USGS:340521117212002:00011:00001",
  "USGS:340521117212003:00011:00001",
  "USGS:11337190:00011:00059",
  "USGS:11337190:00011:00005",
  "USGS:11337190:00011:00060",
  "USGS:11342000:00011:00002",
  "USGS:11342000:00011:00003",
  "USGS:11345500:00011:00001",
  "USGS:11345500:00011:00002",
  "USGS:11348500:00011:00002",
  "USGS:11348500:00011:00003",
  "USGS:11355010:00011:00001",
  "USGS:11355010:00011:00002",
  "USGS:11361000:00011:00001",
  "USGS:11361000:00011:00002",
  "USGS:11370500:00011:00002",
  "USGS:11370500:00011:00003",
  "USGS:11372000:00011:00002",
  "USGS:11372000:00011:00003",
  "USGS:11374000:00011:00002",
  "USGS:11374000:00011:00003",
  "USGS:11376000:00011:00002",
  "USGS:11376000:00011:00003",
  "USGS:11376550:00011:00002",
  "USGS:11376550:00011:00003",
  "USGS:11377100:00011:00002",
  "USGS:11377100:00011:00003",
  "USGS:11379500:00011:00002",
  "USGS:11379500:00011:00003",
  "USGS:11381500:00011:00003",
  "USGS:11381500:00011:00001",
  "USGS:11381500:00011:00002",
  "USGS:11383500:00011:00003",
  "USGS:11383500:00011:00001",
  "USGS:11383500:00011:00002",
  "USGS:11389500:00011:00002",
  "USGS:11389500:00011:00003",
  "USGS:11390000:00011:00001",
  "USGS:11390000:00011:00002",
  "USGS:11390000:00011:00003",
  "USGS:11390500:00011:00001",
  "USGS:11390500:00011:00002",
  "USGS:11390500:00011:00003",
  "USGS:11401920:00011:00002",
  "USGS:11401920:00011:00001",
  "USGS:11402000:00011:00001",
  "USGS:11402000:00011:00002",
  "USGS:11413000:00011:00001",
  "USGS:11413000:00011:00002",
  "USGS:11418500:00011:00002",
  "USGS:11418500:00011:00003",
  "USGS:11421000:00011:00003",
  "USGS:11421000:00011:00004",
  "USGS:11424000:00011:00001",
  "USGS:11424000:00011:00002",
  "USGS:11424500:00011:00002",
  "USGS:11425500:00011:00001",
  "USGS:11425500:00011:00002",
  "USGS:11425500:00011:00003",
  "USGS:11425500:00011:00018",
  "USGS:11425500:00011:00019",
  "USGS:11427000:00011:00002",
  "USGS:11427000:00011:00003",
  "USGS:11433790:00011:00001",
  "USGS:11446030:00011:00001",
  "USGS:11446220:00011:00001",
  "USGS:11446500:00011:00001",
  "USGS:11446500:00011:00002",
  "USGS:11446500:00011:00003",
  "USGS:11446700:00011:00001",
  "USGS:11446980:00011:00001",
  "USGS:11447360:00011:00001",
  "USGS:11447360:00011:00002",
  "USGS:11447650:00011:00001",
  "USGS:11447650:00011:00041",
  "USGS:11447650:00011:00013",
  "USGS:11447650:00011:00002",
  "USGS:11447650:00011:00012",
  "USGS:11447650:00011:00003",
  "USGS:11447650:00011:00047",
  "USGS:11447650:00011:00038",
  "USGS:11447650:00011:00052",
  "USGS:11447650:00011:00009",
  "USGS:11447650:00011:00007",
  "USGS:11447650:00011:00048",
  "USGS:11447650:00011:00050",
  "USGS:11447650:00011:00039",
  "USGS:11447650:00011:00045",
  "USGS:11447650:00011:00011",
  "USGS:11447650:00011:00040",
  "USGS:11447650:00011:00046",
  "USGS:11447830:00011:00008",
  "USGS:11447830:00011:00012",
  "USGS:11447830:00011:00004",
  "USGS:11447830:00011:00011",
  "USGS:11447830:00011:00009",
  "USGS:11447830:00011:00019",
  "USGS:11447830:00011:00020",
  "USGS:11447830:00011:00021",
  "USGS:11447830:00011:00024",
  "USGS:11447830:00011:00015",
  "USGS:11447850:00011:00017",
  "USGS:11447850:00011:00012",
  "USGS:11447850:00011:00001",
  "USGS:11447850:00011:00011",
  "USGS:11447850:00011:00018",
  "USGS:11447850:00011:00019",
  "USGS:11447850:00011:00020",
  "USGS:11447850:00011:00022",
  "USGS:11447850:00011:00024",
  "USGS:11447850:00011:00002",
  "USGS:11447890:00011:00017",
  "USGS:11447890:00011:00012",
  "USGS:11447890:00011:00003",
  "USGS:11447890:00011:00011",
  "USGS:11447890:00011:00019",
  "USGS:11447890:00011:00027",
  "USGS:11447890:00011:00028",
  "USGS:11447890:00011:00020",
  "USGS:11447890:00011:00023",
  "USGS:11447890:00011:00025",
  "USGS:11447890:00011:00024",
  "USGS:11447890:00011:00005",
  "USGS:11447890:00011:00029",
  "USGS:11447903:00011:00012",
  "USGS:11447903:00011:00001",
  "USGS:11447903:00011:00011",
  "USGS:11447903:00011:00024",
  "USGS:11447903:00011:00015",
  "USGS:11447903:00011:00008",
  "USGS:11447905:00011:00012",
  "USGS:11447905:00011:00003",
  "USGS:11447905:00011:00011",
  "USGS:11447905:00011:00004",
  "USGS:11449500:00011:00001",
  "USGS:11449500:00011:00002",
  "USGS:11450000:00011:00002",
  "USGS:11451000:00011:00001",
  "USGS:11451000:00011:00002",
  "USGS:11451100:00011:00001",
  "USGS:11451100:00011:00002",
  "USGS:11451290:00011:00002",
  "USGS:11451290:00011:00001",
  "USGS:11451292:00011:00001",
  "USGS:11451292:00011:00002",
  "USGS:11451292:00011:00013",
  "USGS:11451300:00011:00001",
  "USGS:11451300:00011:00002",
  "USGS:11451715:00011:00002",
  "USGS:11451715:00011:00001",
  "USGS:11452500:00011:00002",
  "USGS:11452500:00011:00003",
  "USGS:02043433:00011:00001",
  "USGS:0204382800:00011:00015",
  "USGS:11133000:00011:00009",
  "USGS:11134000:00011:00001",
  "USGS:11134000:00011:00002",
  "USGS:11135800:00011:00001",
  "USGS:11135800:00011:00002",
  "USGS:11136600:00011:00002",
  "USGS:11136600:00011:00001",
  "USGS:11136800:00011:00001",
  "USGS:11136800:00011:00002",
  "USGS:11137900:00011:00001",
  "USGS:11137900:00011:00002",
  "USGS:11138500:00011:00001",
  "USGS:11138500:00011:00002",
  "USGS:11140000:00011:00005",
  "USGS:11140000:00011:00006",
  "USGS:11140585:00011:00001",
  "USGS:11140585:00011:00002",
  "USGS:11141280:00011:00002",
  "USGS:11141280:00011:00005",
  "USGS:11143000:00011:00002",
  "USGS:11143000:00011:00003",
  "USGS:11143200:00011:00001",
  "USGS:11143200:00011:00002",
  "USGS:11143250:00011:00001",
  "USGS:11143250:00011:00004",
  "USGS:11147500:00011:00001",
  "USGS:11147500:00011:00002",
  "USGS:11148500:00011:00002",
  "USGS:11148900:00011:00002",
  "USGS:11148900:00011:00005",
  "USGS:11149400:00011:00001",
  "USGS:11149400:00011:00002",
  "USGS:11149900:00011:00002",
  "USGS:11149900:00011:00005",
  "USGS:11150500:00011:00001",
  "USGS:11150500:00011:00002",
  "USGS:11151700:00011:00001",
  "USGS:11151700:00011:00002",
  "USGS:11151870:00011:00005",
  "USGS:11152000:00011:00001",
  "USGS:11152000:00011:00002",
  "USGS:11152050:00011:00002",
  "USGS:11152050:00011:00001",
  "USGS:11152300:00011:00002",
  "USGS:11152300:00011:00006",
  "USGS:11152500:00011:00002",
  "USGS:11152500:00011:00006",
  "USGS:11152650:00011:00001",
  "USGS:11152650:00011:00002",
  "USGS:11153000:00011:00001",
  "USGS:11153000:00011:00002",
  "USGS:11153650:00011:00001",
  "USGS:11153650:00011:00002",
  "USGS:11154700:00011:00002",
  "USGS:11154700:00011:00001",
  "USGS:11156500:00011:00001",
  "USGS:11156500:00011:00002",
  "USGS:11157500:00011:00001",
  "USGS:11157500:00011:00002",
  "USGS:11158600:00011:00001",
  "USGS:11158600:00011:00002",
  "USGS:11159000:00011:00002",
  "USGS:11159000:00011:00004",
  "USGS:11159200:00011:00001",
  "USGS:11159200:00011:00002",
  "USGS:11160000:00011:00002",
  "USGS:11160000:00011:00003",
  "USGS:11160500:00011:00002",
  "USGS:11160500:00011:00005",
  "USGS:11161000:00011:00001",
  "USGS:11161000:00011:00002",
  "USGS:11162500:00011:00002",
  "USGS:11162500:00011:00005",
  "USGS:11162570:00011:00001",
  "USGS:11162570:00011:00002",
  "USGS:11162618:00011:00001",
  "USGS:11162620:00011:00013",
  "USGS:11162620:00011:00002",
  "USGS:11162620:00011:00001",
  "USGS:11162630:00011:00001",
  "USGS:11162630:00011:00002",
  "USGS:11162750:00011:00001",
  "USGS:11162753:00011:00003",
  "USGS:11162753:00011:00001",
  "USGS:11162753:00011:00002",
  "USGS:11162765:00011:00001",
  "USGS:11162765:00011:00003",
  "USGS:11162765:00011:00002",
  "USGS:11162765:00011:00004",
  "USGS:11162765:00011:00019",
  "USGS:11480390:00011:00001",
  "USGS:11480390:00011:00002",
  "USGS:11455139:00011:00009",
  "USGS:11455139:00011:00010",
  "USGS:11455139:00011:00004",
  "USGS:11455139:00011:00005",
  "USGS:11455139:00011:00007",
  "USGS:11455139:00011:00006",
  "USGS:11455139:00011:00011",
  "USGS:11455146:00011:00002",
  "USGS:11455146:00011:00003",
  "USGS:11455146:00011:00008",
  "USGS:11455146:00011:00009",
  "USGS:11455146:00011:00004",
  "USGS:11455146:00011:00005",
  "USGS:11455146:00011:00006",
  "USGS:11455146:00011:00010",
  "USGS:11455146:00011:00012",
  "USGS:11455146:00011:00011",
  "USGS:11455146:00011:00001",
  "USGS:11455165:00011:00012",
  "USGS:11455165:00011:00005",
  "USGS:11455165:00011:00011",
  "USGS:11455165:00011:00022",
  "USGS:11455165:00011:00017",
  "USGS:11455165:00011:00015",
  "USGS:11455165:00011:00019",
  "USGS:11455315:00011:00058",
  "USGS:11455315:00011:00003",
  "USGS:11455315:00011:00001",
  "USGS:11455315:00011:00002",
  "USGS:11455315:00011:00059",
  "USGS:11455315:00011:00024",
  "USGS:11455315:00011:00065",
  "USGS:11455315:00011:00066",
  "USGS:11455315:00011:00060",
  "USGS:11455315:00011:00061",
  "USGS:11455315:00011:00069",
  "USGS:11455315:00011:00063",
  "USGS:11455315:00011:00020",
  "USGS:11455315:00011:00062",
  "USGS:11455315:00011:00004",
  "USGS:11455315:00011:00057",
  "USGS:11455315:00011:00022",
  "USGS:11455335:00011:00003",
  "USGS:11455335:00011:00004",
  "USGS:11455335:00011:00002",
  "USGS:11455335:00011:00018",
  "USGS:11455335:00011:00020",
  "USGS:11455335:00011:00005",
  "USGS:11455335:00011:00024",
  "USGS:11455350:00011:00028",
  "USGS:11455350:00011:00012",
  "USGS:11455350:00011:00009",
  "USGS:11455350:00011:00011",
  "USGS:11455350:00011:00029",
  "USGS:11455350:00011:00035",
  "USGS:11455350:00011:00039",
  "USGS:11455350:00011:00030",
  "USGS:11455350:00011:00033",
  "USGS:11455350:00011:00031",
  "USGS:11455350:00011:00022",
  "USGS:11455350:00011:00032",
  "USGS:11455350:00011:00015",
  "USGS:11455350:00011:00036",
  "USGS:11455350:00011:00038",
  "USGS:11455420:00011:00012",
  "USGS:11455420:00011:00005",
  "USGS:11455420:00011:00011",
  "USGS:11455420:00011:00035",
  "USGS:11455420:00011:00006",
  "USGS:11455420:00011:00009",
  "USGS:11455478:00011:00024",
  "USGS:11455478:00011:00002",
  "USGS:11455478:00011:00001",
  "USGS:11455478:00011:00025",
  "USGS:11455478:00011:00058",
  "USGS:11455478:00011:00026",
  "USGS:11455478:00011:00029",
  "USGS:11455478:00011:00027",
  "USGS:11455478:00011:00028",
  "USGS:11455478:00011:00059",
  "USGS:11455780:00011:00005",
  "USGS:11455780:00011:00006",
  "USGS:11455780:00011:00003",
  "USGS:11455780:00011:00004",
  "USGS:11455780:00011:00015",
  "USGS:11455780:00011:00009",
  "USGS:11461500:00011:00005",
  "USGS:11455780:00011:00010",
  "USGS:11455780:00011:00007",
  "USGS:11455780:00011:00008",
  "USGS:11456000:00011:00002",
  "USGS:11456000:00011:00005",
  "USGS:11458000:00011:00002",
  "USGS:11458000:00011:00006",
  "USGS:11458433:00011:00003",
  "USGS:11458433:00011:00002",
  "USGS:11458433:00011:00001",
  "USGS:11458433:00011:00004",
  "USGS:11458500:00011:00001",
  "USGS:11458500:00011:00002",
  "USGS:11459150:00011:00003",
  "USGS:11459150:00011:00001",
  "USGS:11459150:00011:00005",
  "USGS:11459500:00011:00001",
  "USGS:11459500:00011:00002",
  "USGS:11460000:00011:00002",
  "USGS:11460000:00011:00005",
  "USGS:11460151:00011:00002",
  "USGS:11460400:00011:00001",
  "USGS:11460400:00011:00002",
  "USGS:11460600:00011:00001",
  "USGS:11460600:00011:00002",
  "USGS:11460750:00011:00001",
  "USGS:11460750:00011:00002",
  "USGS:11461000:00011:00002",
  "USGS:11461000:00011:00005",
  "USGS:11461500:00011:00002",
  "USGS:11462080:00011:00002",
  "USGS:11462080:00011:00001",
  "USGS:11462500:00011:00001",
  "USGS:11462500:00011:00002",
  "USGS:11462500:00011:00003",
  "USGS:11462500:00011:00015",
  "USGS:11462500:00011:00016",
  "USGS:11462500:00011:00017",
  "USGS:11462500:00011:00021",
  "USGS:11463000:00011:00003",
  "USGS:11463000:00011:00004",
  "USGS:11463000:00011:00007",
  "USGS:11463000:00011:00002",
  "USGS:11463170:00011:00001",
  "USGS:11463170:00011:00002",
  "USGS:11463200:00011:00002",
  "USGS:11463200:00011:00005",
  "USGS:11463500:00011:00001",
  "USGS:11463500:00011:00002",
  "USGS:11463682:00011:00003",
  "USGS:11463682:00011:00002",
  "USGS:11463682:00011:00001",
  "USGS:11463682:00011:00005",
  "USGS:11463682:00011:00004",
  "USGS:11463682:00011:00015",
  "USGS:11463682:00011:00016",
  "USGS:11463900:00011:00001",
  "USGS:11463900:00011:00002",
  "USGS:11463980:00011:00003",
  "USGS:11463980:00011:00002",
  "USGS:11463980:00011:00001",
  "USGS:11463980:00011:00004",
  "USGS:11463980:00011:00005",
  "USGS:11463980:00011:00007",
  "USGS:11463980:00011:00011",
  "USGS:11464000:00011:00002",
  "USGS:11464000:00011:00003",
  "USGS:11465200:00011:00002",
  "USGS:11465200:00011:00005",
  "USGS:11465240:00011:00003",
  "USGS:11465240:00011:00002",
  "USGS:11465240:00011:00001",
  "USGS:11465240:00011:00004",
  "USGS:11465240:00011:00005",
  "USGS:11465240:00011:00006",
  "USGS:11465240:00011:00007",
  "USGS:11465240:00011:00090",
  "USGS:11465240:00011:00091",
  "USGS:11465350:00011:00001",
  "USGS:11465350:00011:00002",
  "USGS:11465390:00011:00003",
  "USGS:11465390:00011:00001",
  "USGS:11465660:00011:00002",
  "USGS:11465660:00011:00001",
  "USGS:11465680:00011:00001",
  "USGS:11465680:00011:00002",
  "USGS:11465690:00011:00002",
  "USGS:11465690:00011:00001",
  "USGS:11465700:00011:00001",
  "USGS:11465700:00011:00002",
  "USGS:11465750:00011:00002",
  "USGS:11465750:00011:00001",
  "USGS:11466170:00011:00004",
  "USGS:11466170:00011:00002",
  "USGS:11466200:00011:00001",
  "USGS:11466200:00011:00002",
  "USGS:08355050:00011:00010",
  "USGS:08355050:00011:00011",
  "USGS:08355490:00011:00001",
  "USGS:08355490:00011:00002",
  "USGS:08358300:00011:00006",
  "USGS:08358300:00011:00010",
  "USGS:08358400:00011:00005",
  "USGS:08358400:00011:00009",
  "USGS:08359500:00011:00001",
  "USGS:08359500:00011:00002",
  "USGS:08361000:00011:00004",
  "USGS:08361000:00011:00005",
  "USGS:08377900:00011:00006",
  "USGS:08377900:00011:00001",
  "USGS:08377900:00011:00002",
  "USGS:08378500:00011:00005",
  "USGS:08378500:00011:00006",
  "USGS:08379500:00011:00001",
  "USGS:08379500:00011:00002",
  "USGS:08380500:00011:00001",
  "USGS:08380500:00011:00002",
  "USGS:08382500:00011:00001",
  "USGS:08382500:00011:00002",
  "USGS:08382600:00011:00004",
  "USGS:08382600:00011:00005",
  "USGS:08382650:00011:00004",
  "USGS:11276500:00011:00003",
  "USGS:11276600:00011:00001",
  "USGS:11276600:00011:00002",
  "USGS:11276600:00011:00003",
  "USGS:11276900:00011:00003",
  "USGS:11276900:00011:00001",
  "USGS:11276900:00011:00002",
  "USGS:11277100:00011:00001",
  "USGS:11277200:00011:00001",
  "USGS:11277200:00011:00003",
  "USGS:11277300:00011:00014",
  "USGS:11277300:00011:00001",
  "USGS:11277300:00011:00002",
  "USGS:11277500:00011:00001",
  "USGS:11277500:00011:00002",
  "USGS:11278000:00011:00001",
  "USGS:11278000:00011:00004",
  "USGS:11278000:00011:00005",
  "USGS:11278300:00011:00003",
  "USGS:11278300:00011:00001",
  "USGS:11278300:00011:00002",
  "USGS:11278400:00011:00003",
  "USGS:11278400:00011:00001",
  "USGS:11278400:00011:00002",
  "USGS:11284400:00011:00001",
  "USGS:11284400:00011:00002",
  "USGS:11285500:00011:00003",
  "USGS:11285500:00011:00001",
  "USGS:11285500:00011:00002",
  "USGS:11285500:00011:00004",
  "USGS:11285500:00011:00006",
  "USGS:11285500:00011:00007",
  "USGS:11285500:00011:00005",
  "USGS:11287500:00011:00001",
  "USGS:11287500:00011:00002",
  "USGS:11289000:00011:00001",
  "USGS:11289000:00011:00002",
  "USGS:11289500:00011:00001",
  "USGS:11289650:00011:00001",
  "USGS:11289650:00011:00002",
  "USGS:11289650:00011:00003",
  "USGS:11290000:00011:00001",
  "USGS:11290000:00011:00002",
  "USGS:11290000:00011:00003",
  "USGS:11290000:00011:00004",
  "USGS:11299600:00011:00001",
  "USGS:11299600:00011:00002",
  "USGS:11302000:00011:00001",
  "USGS:11302500:00011:00001",
  "USGS:11303000:00011:00001",
  "USGS:11303000:00011:00002",
  "USGS:11303000:00011:00003",
  "USGS:11303000:00011:00004",
  "USGS:11303500:00011:00003",
  "USGS:11303500:00011:00004",
  "USGS:11303500:00011:00005",
  "USGS:11304810:00011:00012",
  "USGS:11304810:00011:00005",
  "USGS:11304810:00011:00011",
  "USGS:11304810:00011:00024",
  "USGS:11304810:00011:00006",
  "USGS:11304810:00011:00030",
  "USGS:11311300:00011:00012",
  "USGS:11311300:00011:00001",
  "USGS:11311300:00011:00011",
  "USGS:11311300:00011:00002",
  "USGS:11312672:00011:00012",
  "USGS:11312672:00011:00001",
  "USGS:11312672:00011:00011",
  "USGS:11312672:00011:00002",
  "USGS:11312676:00011:00012",
  "USGS:11312676:00011:00002",
  "USGS:11312676:00011:00011",
  "USGS:11312676:00011:00025",
  "USGS:11312676:00011:00005",
  "USGS:11312676:00011:00029",
  "USGS:11312685:00011:00003",
  "USGS:11312685:00011:00004",
  "USGS:11312685:00011:00002",
  "USGS:11312685:00011:00005",
  "USGS:11312968:00011:00012",
  "USGS:11312968:00011:00003",
  "USGS:11312968:00011:00011",
  "USGS:11312968:00011:00004",
  "USGS:11313240:00011:00012",
  "USGS:11313240:00011:00003",
  "USGS:11313240:00011:00004",
  "USGS:11313315:00011:00012",
  "USGS:11313315:00011:00003",
  "USGS:11313315:00011:00011",
  "USGS:11313315:00011:00004",
  "USGS:11313405:00011:00012",
  "USGS:11313405:00011:00002",
  "USGS:11313405:00011:00011",
  "USGS:11313405:00011:00005",
  "USGS:11313405:00011:00029",
  "USGS:11313431:00011:00003",
  "USGS:11313431:00011:00004",
  "USGS:11313431:00011:00002",
  "USGS:11313431:00011:00005",
  "USGS:11313433:00011:00022",
  "USGS:11313433:00011:00012",
  "USGS:11313433:00011:00005",
  "USGS:11313433:00011:00023",
  "USGS:11313433:00011:00001",
  "USGS:11313433:00011:00027",
  "USGS:11313433:00011:00006",
  "USGS:11313434:00011:00003",
  "USGS:11313434:00011:00004",
  "USGS:11313434:00011:00002",
  "USGS:11313434:00011:00005",
  "USGS:11313440:00011:00003",
  "USGS:11313440:00011:00004",
  "USGS:11313440:00011:00002",
  "USGS:11313440:00011:00005",
  "USGS:11313452:00011:00003",
  "USGS:11313452:00011:00004",
  "USGS:11313452:00011:00002",
  "USGS:11313452:00011:00005",
  "USGS:11313460:00011:00003",
  "USGS:11313460:00011:00004",
  "USGS:11313460:00011:00002",
  "USGS:11313460:00011:00005",
  "USGS:11335000:00011:00001",
  "USGS:11335000:00011:00002",
  "USGS:11335000:00011:00003",
  "USGS:11336580:00011:00001",
  "USGS:11336580:00011:00002",
  "USGS:11336585:00011:00002",
  "USGS:11336585:00011:00001",
  "USGS:11336600:00011:00012",
  "USGS:11336600:00011:00006",
  "USGS:11336600:00011:00011",
  "USGS:11336600:00011:00001",
  "USGS:11336680:00011:00003",
  "USGS:11336680:00011:00001",
  "USGS:11336680:00011:00002",
  "USGS:11336680:00011:00020",
  "USGS:11336680:00011:00004",
  "USGS:11336680:00011:00022",
  "USGS:11336685:00011:00003",
  "USGS:11336685:00011:00001",
  "USGS:11336685:00011:00020",
  "USGS:11336685:00011:00004",
  "USGS:11336685:00011:00022",
  "USGS:11336790:00011:00003",
  "USGS:11336790:00011:00004",
  "USGS:11336790:00011:00002",
  "USGS:11336790:00011:00014",
  "USGS:11336790:00011:00005",
  "USGS:11336790:00011:00016",
  "USGS:07047855:00011:00003",
  "USGS:07047855:00011:00004",
  "USGS:07047855:00011:00002",
  "USGS:07047855:00011:00014",
  "USGS:07047855:00011:00001",
  "USGS:11469000:00011:00002",
  "USGS:11469000:00011:00003",
  "USGS:11473900:00011:00003",
  "USGS:11473900:00011:00007",
  "USGS:11475000:00011:00002",
  "USGS:11475000:00011:00005",
  "USGS:11475560:00011:00001",
  "USGS:11475560:00011:00002",
  "USGS:11475560:00011:00005",
  "USGS:11475610:00011:00003",
  "USGS:11475610:00011:00002",
  "USGS:11475610:00011:00001",
  "USGS:11475800:00011:00002",
  "USGS:11475800:00011:00003",
  "USGS:11476500:00011:00002",
  "USGS:11476500:00011:00005",
  "USGS:11476600:00011:00002",
  "USGS:11476600:00011:00005",
  "USGS:11477000:00011:00002",
  "USGS:11477000:00011:00006",
  "USGS:11478500:00011:00002",
  "USGS:11478500:00011:00003",
  "USGS:11479560:00011:00001",
  "USGS:11481000:00011:00002",
  "USGS:11481000:00011:00005",
  "USGS:11481200:00011:00001",
  "USGS:11481200:00011:00002",
  "USGS:11481500:00011:00002",
  "USGS:11481500:00011:00005",
  "USGS:11482500:00011:00002",
  "USGS:11482500:00011:00005",
  "USGS:11516530:00011:00004",
  "USGS:11516530:00011:00005",
  "USGS:11517000:00011:00001",
  "USGS:11517000:00011:00002",
  "USGS:11517500:00011:00002",
  "USGS:11517500:00011:00003",
  "USGS:11519500:00011:00002",
  "USGS:11519500:00011:00003",
  "USGS:11520500:00011:00002",
  "USGS:11520500:00011:00003",
  "USGS:11521500:00011:00001",
  "USGS:11521500:00011:00002",
  "USGS:11522500:00011:00004",
  "USGS:11522500:00011:00005",
  "USGS:11523000:00011:00001",
  "USGS:11523000:00011:00002",
  "USGS:11523000:00011:00005",
  "USGS:11523200:00011:00001",
  "USGS:11523200:00011:00002",
  "USGS:11525500:00011:00002",
  "USGS:11525500:00011:00003",
  "USGS:11525530:00011:00001",
  "USGS:11525530:00011:00002",
  "USGS:11525630:00011:00001",
  "USGS:11525630:00011:00002",
  "USGS:11525655:00011:00002",
  "USGS:11525655:00011:00005",
  "USGS:11525670:00011:00001",
  "USGS:11525670:00011:00002",
  "USGS:11525854:00011:00001",
  "USGS:11525854:00011:00002",
  "USGS:11526250:00011:00001",
  "USGS:11526250:00011:00002",
  "USGS:11526400:00011:00001",
  "USGS:11526400:00011:00002",
  "USGS:11526500:00011:00002",
  "USGS:11526500:00011:00005",
  "USGS:11527000:00011:00002",
  "USGS:11527000:00011:00003",
  "USGS:11528700:00011:00002",
  "USGS:11528700:00011:00005",
  "USGS:11530000:00011:00001",
  "USGS:11530000:00011:00002",
  "USGS:11530000:00011:00005",
  "USGS:11530500:00011:00006",
  "USGS:11530500:00011:00002",
  "USGS:11530500:00011:00004",
  "USGS:11532500:00011:00002",
  "USGS:11532500:00011:00006",
  "USGS:11532650:00011:00001",
  "USGS:323313117033901:00011:00001",
  "USGS:07048490:00011:00013",
  "USGS:07048490:00011:00002",
  "USGS:07048490:00011:00003",
  "USGS:07048490:00011:00001",
  "USGS:07048550:00011:00017",
  "USGS:07048550:00011:00012",
  "USGS:07048550:00011:00001",
  "USGS:07048550:00011:00018",
  "USGS:07048550:00011:00019",
  "USGS:07048600:00011:00005",
  "USGS:07048600:00011:00004",
  "USGS:323527117050001:00011:00001",
  "USGS:323527117050002:00011:00001",
  "USGS:323527117050003:00011:00001",
  "USGS:323527117050004:00011:00001",
  "USGS:323527117050005:00011:00001",
  "USGS:323528117031401:00011:00001",
  "USGS:323528117031402:00011:00001",
  "USGS:323528117031403:00011:00001",
  "USGS:323528117031404:00011:00001",
  "USGS:323528117031405:00011:00001",
  "USGS:323659117033301:00011:00001",
  "USGS:323659117033302:00011:00001",
  "USGS:323659117033303:00011:00001",
  "USGS:323659117033304:00011:00001",
  "USGS:323659117033305:00011:00001",
  "USGS:323659117033306:00011:00001",
  "USGS:323908116512401:00011:00001",
  "USGS:323915117055301:00011:00001",
  "USGS:323915117055302:00011:00001",
  "USGS:323915117055303:00011:00001",
  "USGS:323915117055304:00011:00001",
  "USGS:323915117055305:00011:00001",
  "USGS:323932117050801:00011:00090",
  "USGS:323932117050801:00011:00001",
  "USGS:323932117050802:00011:00002",
  "USGS:323932117050802:00011:00001",
  "USGS:323932117050803:00011:00001",
  "USGS:323932117050804:00011:00001",
  "USGS:323932117050805:00011:00001",
  "USGS:323932117050806:00011:00001",
  "USGS:324055117064401:00011:00001",
  "USGS:324055117064402:00011:00001",
  "USGS:324055117064403:00011:00001",
  "USGS:324055117064404:00011:00001",
  "USGS:324055117064405:00011:00001",
  "USGS:324116117050801:00011:00001",
  "USGS:324116117050802:00011:00001",
  "USGS:324116117050803:00011:00001",
  "USGS:324116117050804:00011:00001",
  "USGS:324116117050805:00011:00001",
  "USGS:324307117063501:00011:00001",
  "USGS:324307117063502:00011:00001",
  "USGS:324307117063503:00011:00001",
  "USGS:324307117063504:00011:00001",
  "USGS:324307117063505:00011:00001",
  "USGS:324307117063506:00011:00001",
  "USGS:324318117083101:00011:00001",
  "USGS:324318117083102:00011:00001",
  "USGS:07358550:00011:00002",
  "USGS:07358550:00011:00003",
  "USGS:07358550:00011:00004",
  "USGS:07358550:00011:00001",
  "USGS:07358570:00011:00004",
  "USGS:07358570:00011:00001",
  "USGS:07359002:00011:00003",
  "USGS:07359002:00011:00013",
  "USGS:07359002:00011:00002",
  "USGS:07359002:00011:00001",
  "USGS:07359610:00011:00022",
  "USGS:07359610:00011:00002",
  "USGS:07359610:00011:00001",
  "USGS:07360200:00011:00012",
  "USGS:330514116582901:00011:00001",
  "USGS:330514116582902:00011:00001",
  "USGS:330514116582903:00011:00001",
  "USGS:330555117010101:00011:00002",
  "USGS:330555117010101:00011:00001",
  "USGS:330555117010102:00011:00002",
  "USGS:330555117010102:00011:00001",
  "USGS:330555117010103:00011:00002",
  "USGS:330555117010103:00011:00001",
  "USGS:332535117341001:00011:00001",
  "USGS:332747117061101:00011:00001",
  "USGS:332747117061102:00011:00001",
  "USGS:332819117070601:00011:00001",
  "USGS:332819117070602:00011:00001",
  "USGS:332819117070603:00011:00001",
  "USGS:332819117070604:00011:00001",
  "USGS:332819117070605:00011:00001",
  "USGS:332819117070606:00011:00001",
  "USGS:332857117043301:00011:00001",
  "USGS:332857117043302:00011:00001",
  "USGS:332857117043303:00011:00001",
  "USGS:332857117043304:00011:00001",
  "USGS:332857117043305:00011:00001",
  "USGS:332944116583301:00011:00003",
  "USGS:333001117005701:00011:00001",
  "USGS:333001117005702:00011:00001",
  "USGS:333001117005703:00011:00001",
  "USGS:333001117005705:00011:00001",
  "USGS:340046117020801:00011:00001",
  "USGS:340046117020802:00011:00001",
  "USGS:340046117020803:00011:00001",
  "USGS:340046117020804:00011:00001",
  "USGS:340130117054901:00011:00001",
  "USGS:340130117054902:00011:00001",
  "USGS:340130117054903:00011:00001",
  "USGS:340130117054904:00011:00001",
  "USGS:07075270:00011:00004",
  "USGS:07075270:00011:00002",
  "USGS:07075270:00011:00007",
  "USGS:07075270:00011:00001",
  "USGS:07075270:00011:00005",
  "USGS:07075270:00011:00006",
  "USGS:07075270:00011:00008",
  "USGS:07075270:00011:00009",
  "USGS:07075270:00011:00010",
  "USGS:07075300:00011:00004",
  "USGS:07075300:00011:00002",
  "USGS:07075300:00011:00003",
  "USGS:07076000:00011:00001",
  "USGS:07076000:00011:00005",
  "USGS:07076506:00011:00004",
  "USGS:07076506:00011:00005",
  "USGS:07076506:00011:00003",
  "USGS:07076506:00011:00001",
  "USGS:07076517:00011:00002",
  "USGS:07076517:00011:00001",
  "USGS:07076530:00011:00003",
  "USGS:07076530:00011:00001",
  "USGS:07076530:00011:00002",
  "USGS:07076634:00011:00003",
  "USGS:07076634:00011:00002",
  "USGS:02081054:00011:00001",
  "USGS:02081094:00011:00001",
  "USGS:02081094:00011:00003",
  "USGS:02081094:00011:00002",
  "USGS:02081094:00011:00006",
  "USGS:02081094:00011:00005",
  "USGS:02081094:00011:00008",
  "USGS:08271000:00011:00001",
  "USGS:08271000:00011:00002",
  "USGS:08275500:00011:00001",
  "USGS:08275500:00011:00002",
  "USGS:08276300:00011:00001",
  "USGS:08276300:00011:00002",
  "USGS:08276500:00011:00001",
  "USGS:08276500:00011:00002",
  "USGS:08277470:00011:00002",
  "USGS:08277470:00011:00001",
  "USGS:08279000:00011:00001",
  "USGS:08279000:00011:00002",
  "USGS:08279500:00011:00006",
  "USGS:08279500:00011:00007",
  "USGS:08281400:00011:00002",
  "USGS:08282300:00011:00001",
  "USGS:08284100:00011:00001",
  "USGS:08284100:00011:00002",
  "USGS:08285500:00011:00001",
  "USGS:08285500:00011:00002",
  "USGS:08286500:00011:00001",
  "USGS:08286500:00011:00002",
  "USGS:08287000:00011:00005",
  "USGS:08287000:00011:00006",
  "USGS:08289000:00011:00001",
  "USGS:08289000:00011:00002",
  "USGS:08290000:00011:00006",
  "USGS:08290000:00011:00007",
  "USGS:08291000:00011:00001",
  "USGS:08291000:00011:00002",
  "USGS:08294200:00011:00001",
  "USGS:08294200:00011:00002",
  "USGS:08294210:00011:00001",
  "USGS:08294210:00011:00002",
  "USGS:08302500:00011:00001",
  "USGS:08302500:00011:00004",
  "USGS:08313000:00011:00009",
  "USGS:08313000:00011:00013",
  "USGS:08313500:00011:00001",
  "USGS:08313500:00011:00002",
  "USGS:08314000:00011:00001",
  "USGS:08314000:00011:00002",
  "USGS:08315480:00011:00004",
  "USGS:08315480:00011:00003",
  "USGS:08315500:00011:00001",
  "USGS:08315500:00011:00004",
  "USGS:08315500:00011:00002",
  "USGS:08316000:00011:00001",
  "USGS:08316000:00011:00002",
  "USGS:08316500:00011:00001",
  "USGS:08316500:00011:00002",
  "USGS:08317200:00011:00001",
  "USGS:08317200:00011:00002",
  "USGS:08317400:00011:00005",
  "USGS:08317400:00011:00006",
  "USGS:08317400:00011:00010",
  "USGS:08317400:00011:00007",
  "USGS:08317400:00011:00020",
  "USGS:08317400:00011:00021",
  "USGS:08317400:00011:00019",
  "USGS:08317950:00011:00005",
  "USGS:08317950:00011:00006",
  "USGS:08319000:00011:00001",
  "USGS:08319000:00011:00002",
  "USGS:08324000:00011:00005",
  "USGS:08324000:00011:00006",
  "USGS:08328950:00011:00002",
  "USGS:08328950:00011:00001",
  "USGS:08329900:00011:00003",
  "USGS:08329900:00011:00001",
  "USGS:08329900:00011:00002",
  "USGS:08329918:00011:00012",
  "USGS:08329918:00011:00002",
  "USGS:08329918:00011:00001",
  "USGS:08329928:00011:00002",
  "USGS:08329928:00011:00001",
  "USGS:08330000:00011:00003",
  "USGS:08330000:00011:00010",
  "USGS:08330600:00011:00001",
  "USGS:08330600:00011:00002",
  "USGS:08330775:00011:00014",
  "USGS:08330775:00011:00001",
  "USGS:08330775:00011:00002",
  "USGS:08330875:00011:00011",
  "USGS:08330875:00011:00001",
  "USGS:08331160:00011:00002",
  "USGS:08331160:00011:00001",
  "USGS:08331510:00011:00010",
  "USGS:08331510:00011:00011",
  "USGS:08332010:00011:00002",
  "USGS:08332010:00011:00006",
  "USGS:08334000:00011:00005",
  "USGS:08334000:00011:00008",
  "USGS:08340500:00011:00001",
  "USGS:08340500:00011:00004",
  "USGS:08341400:00011:00001",
  "USGS:08341400:00011:00002",
  "USGS:08343500:00011:00001",
  "USGS:08343500:00011:00002",
  "USGS:08353000:00011:00002",
  "USGS:08353000:00011:00006",
  "USGS:08354900:00011:00005",
  "USGS:08354900:00011:00009",
  "USGS:06613950:00011:00003",
  "USGS:06613950:00011:00001",
  "USGS:06613950:00011:00004",
  "USGS:06614800:00011:00001",
  "USGS:06614800:00011:00003",
  "USGS:06620000:00011:00005",
  "USGS:06620000:00011:00018",
  "USGS:06620000:00011:00009",
  "USGS:06696980:00011:00004",
  "USGS:06696980:00011:00005",
  "USGS:340521117212004:00011:00001",
  "USGS:340521117212005:00011:00001",
  "USGS:340541117074401:00011:00001",
  "USGS:340541117074402:00011:00001",
  "USGS:340541117074403:00011:00001",
  "USGS:340541117074404:00011:00001",
  "USGS:340541117074405:00011:00001",
  "USGS:340541117074406:00011:00001",
  "USGS:340615117170902:00011:00001",
  "USGS:340615117170903:00011:00001",
  "USGS:340615117170904:00011:00001",
  "USGS:340655117184004:00011:00001",
  "USGS:340655117184005:00011:00001",
  "USGS:340655117184006:00011:00001",
  "USGS:340707117162706:00011:00002",
  "USGS:340707117162706:00011:00001",
  "USGS:340707117162707:00011:00001",
  "USGS:340707117162708:00011:00001",
  "USGS:340716117230601:00011:00001",
  "USGS:340716117230602:00011:00001",
  "USGS:340716117230603:00011:00001",
  "USGS:340716117230604:00011:00001",
  "USGS:340716117230605:00011:00001",
  "USGS:340742117161701:00011:00001",
  "USGS:340800117235901:00011:00001",
  "USGS:340800117235902:00011:00001",
  "USGS:07260671:00011:00003",
  "USGS:07260671:00011:00001",
  "USGS:072606713:00011:00004",
  "USGS:072606713:00011:00001",
  "USGS:07048600:00011:00002",
  "USGS:07048600:00011:00003",
  "USGS:07048600:00011:00001",
  "USGS:07048600:00011:00020",
  "USGS:07048600:00011:00018",
  "USGS:07048600:00011:00019",
  "USGS:07048800:00011:00002",
  "USGS:07048800:00011:00001",
  "USGS:07049000:00011:00005",
  "USGS:07049000:00011:00002",
  "USGS:07049691:00011:00003",
  "USGS:07049691:00011:00002",
  "USGS:07050500:00011:00004",
  "USGS:07050500:00011:00001",
  "USGS:07050500:00011:00003",
  "USGS:07053207:00011:00001",
  "USGS:07053250:00011:00004",
  "USGS:07053250:00011:00001",
  "USGS:07054410:00011:00012",
  "USGS:07054501:00011:00002",
  "USGS:07054501:00011:00001",
  "USGS:07054502:00011:00002",
  "USGS:07054502:00011:00001",
  "USGS:07054527:00011:00002",
  "USGS:07054527:00011:00001",
  "USGS:07055607:00011:00003",
  "USGS:07055607:00011:00004",
  "USGS:07055607:00011:00002",
  "USGS:07055646:00011:00002",
  "USGS:07055646:00011:00014",
  "USGS:07055646:00011:00003",
  "USGS:07055646:00011:00001",
  "USGS:07055660:00011:00003",
  "USGS:07055660:00011:00015",
  "USGS:07055660:00011:00014",
  "USGS:07055660:00011:00016",
  "USGS:07055660:00011:00004",
  "USGS:07055660:00011:00002",
  "USGS:07055660:00011:00001",
  "USGS:07055680:00011:00003",
  "USGS:07055680:00011:00014",
  "USGS:07055680:00011:00002",
  "USGS:07055680:00011:00001",
  "USGS:07055780:00011:00003",
  "USGS:07055780:00011:00001",
  "USGS:07055790:00011:00005",
  "USGS:07055790:00011:00003",
  "USGS:07055790:00011:00001",
  "USGS:07055790:00011:00006",
  "USGS:07055814:00011:00005",
  "USGS:07055814:00011:00004",
  "USGS:07055814:00011:00001",
  "USGS:07055814:00011:00006",
  "USGS:07055814:00011:00009",
  "USGS:07055814:00011:00007",
  "USGS:07055814:00011:00010",
  "USGS:07055814:00011:00008",
  "USGS:07055875:00011:00011",
  "USGS:07055875:00011:00001",
  "USGS:07056000:00011:00004",
  "USGS:07056000:00011:00002",
  "USGS:07056000:00011:00003",
  "USGS:07056515:00011:00002",
  "USGS:07056515:00011:00018",
  "USGS:07056515:00011:00004",
  "USGS:07056515:00011:00001",
  "USGS:07056515:00011:00030",
  "USGS:07056515:00011:00032",
  "USGS:07056515:00011:00029",
  "USGS:07056515:00011:00028",
  "USGS:07056515:00011:00031",
  "USGS:07056700:00011:00002",
  "USGS:07056700:00011:00003",
  "USGS:07056700:00011:00001",
  "USGS:07057370:00011:00002",
  "USGS:07057370:00011:00001",
  "USGS:07058980:00011:00002",
  "USGS:07058980:00011:00012",
  "USGS:07058980:00011:00001",
  "USGS:07059450:00011:00013",
  "USGS:07059450:00011:00001",
  "USGS:07059998:00011:00002",
  "USGS:07059998:00011:00001",
  "USGS:07059998:00011:00003",
  "USGS:07060000:00011:00015",
  "USGS:07060000:00011:00014",
  "USGS:07060001:00011:00002",
  "USGS:07060001:00011:00001",
  "USGS:07060500:00011:00018",
  "USGS:07060500:00011:00004",
  "USGS:07060500:00011:00002",
  "USGS:07060500:00011:00003",
  "USGS:07060710:00011:00016",
  "USGS:07060710:00011:00006",
  "USGS:07060710:00011:00005",
  "USGS:07060728:00011:00002",
  "USGS:07060728:00011:00001",
  "USGS:07061000:00011:00004",
  "USGS:07061000:00011:00002",
  "USGS:07061000:00011:00003",
  "USGS:07064000:00011:00003",
  "USGS:07064000:00011:00001",
  "USGS:07064000:00011:00002",
  "USGS:07069000:00011:00002",
  "USGS:07069000:00011:00005",
  "USGS:07069000:00011:00001",
  "USGS:07069190:00011:00013",
  "USGS:07069190:00011:00015",
  "USGS:07069190:00011:00014",
  "USGS:07069190:00011:00002",
  "USGS:07069190:00011:00001",
  "USGS:07069220:00011:00015",
  "USGS:07069220:00011:00014",
  "USGS:07069220:00011:00001",
  "USGS:07069295:00011:00004",
  "USGS:07069295:00011:00002",
  "USGS:07069295:00011:00001",
  "USGS:07069305:00011:00002",
  "USGS:07069305:00011:00004",
  "USGS:07069305:00011:00001",
  "USGS:07069500:00011:00004",
  "USGS:07069500:00011:00002",
  "USGS:07069500:00011:00003",
  "USGS:07072000:00011:00004",
  "USGS:07072000:00011:00002",
  "USGS:07072000:00011:00003",
  "USGS:07072500:00011:00001",
  "USGS:07072500:00011:00002",
  "USGS:07074000:00011:00004",
  "USGS:07074000:00011:00003",
  "USGS:07074420:00011:00002",
  "USGS:07074420:00011:00003",
  "USGS:07074420:00011:00001",
  "USGS:07074500:00011:00004",
  "USGS:07074500:00011:00002",
  "USGS:07074500:00011:00003",
  "USGS:07074850:00011:00014",
  "USGS:07074850:00011:00002",
  "USGS:07075000:00011:00003",
  "USGS:07075000:00011:00005",
  "USGS:07075000:00011:00002",
  "USGS:07075250:00011:00005",
  "USGS:07075250:00011:00002",
  "USGS:07075250:00011:00021",
  "USGS:07075250:00011:00001",
  "USGS:07075250:00011:00006",
  "USGS:07075250:00011:00007",
  "USGS:07075250:00011:00008",
  "USGS:07075250:00011:00009",
  "USGS:07075250:00011:00023",
  "USGS:343056093030901:00011:00001",
  "USGS:06713500:00011:00001",
  "USGS:06713500:00011:00002",
  "USGS:06714215:00011:00001",
  "USGS:06714215:00011:00006",
  "USGS:06714360:00011:00002",
  "USGS:08382650:00011:00005",
  "USGS:08382830:00011:00004",
  "USGS:08382830:00011:00005",
  "USGS:08383500:00011:00001",
  "USGS:08383500:00011:00002",
  "USGS:08384500:00011:00001",
  "USGS:08384500:00011:00002",
  "USGS:08385000:00011:00001",
  "USGS:08385000:00011:00002",
  "USGS:08385503:00011:00002",
  "USGS:08385503:00011:00001",
  "USGS:08385522:00011:00002",
  "USGS:08385522:00011:00001",
  "USGS:08385630:00011:00002",
  "USGS:08385630:00011:00001",
  "USGS:08386000:00011:00004",
  "USGS:08386000:00011:00016",
  "USGS:08386505:00011:00002",
  "USGS:08386505:00011:00001",
  "USGS:08387000:00011:00001",
  "USGS:08387000:00011:00002",
  "USGS:08387550:00011:00014",
  "USGS:08387550:00011:00013",
  "USGS:08387575:00011:00002",
  "USGS:08387575:00011:00001",
  "USGS:08387600:00011:00001",
  "USGS:08387600:00011:00002",
  "USGS:08388450:00011:00004",
  "USGS:08388450:00011:00001",
  "USGS:08388500:00011:00001",
  "USGS:08390020:00011:00002",
  "USGS:08390020:00011:00001",
  "USGS:08390500:00011:00004",
  "USGS:08390500:00011:00005",
  "USGS:08390800:00011:00004",
  "USGS:08390800:00011:00005",
  "USGS:08393610:00011:00002",
  "USGS:08393610:00011:00001",
  "USGS:08394024:00011:00002",
  "USGS:08394024:00011:00001",
  "USGS:08394033:00011:00002",
  "USGS:08394033:00011:00001",
  "USGS:08394500:00011:00001",
  "USGS:08394500:00011:00002",
  "USGS:08395500:00011:00001",
  "USGS:08395500:00011:00002",
  "USGS:08396500:00011:00005",
  "USGS:08396500:00011:00021",
  "USGS:08397600:00011:00001",
  "USGS:08397600:00011:00002",
  "USGS:08397620:00011:00002",
  "USGS:08397620:00011:00001",
  "USGS:08398500:00011:00001",
  "USGS:08398500:00011:00002",
  "USGS:08399500:00011:00001",
  "USGS:08399500:00011:00002",
  "USGS:08400000:00011:00001",
  "USGS:08400000:00011:00002",
  "USGS:08401200:00011:00001",
  "USGS:08401200:00011:00002",
  "USGS:08401500:00011:00001",
  "USGS:08401500:00011:00002",
  "USGS:08401900:00011:00001",
  "USGS:08401900:00011:00002",
  "USGS:08402000:00011:00005",
  "USGS:08402000:00011:00006",
  "USGS:08403500:00011:00001",
  "USGS:08403500:00011:00002",
  "USGS:08404000:00011:00001",
  "USGS:08404000:00011:00002",
  "USGS:08405105:00011:00002",
  "USGS:08405105:00011:00001",
  "USGS:08405150:00011:00001",
  "USGS:08405150:00011:00002",
  "USGS:07103755:00011:00001",
  "USGS:07103755:00011:00002",
  "USGS:07103780:00011:00001",
  "USGS:07103780:00011:00003",
  "USGS:07103797:00011:00002",
  "USGS:07103797:00011:00006",
  "USGS:07103800:00011:00013",
  "USGS:07103800:00011:00001",
  "USGS:07103800:00011:00003",
  "USGS:07103970:00011:00017",
  "USGS:07103970:00011:00002",
  "USGS:07103970:00011:00001",
  "USGS:07103970:00011:00014",
  "USGS:07103970:00011:00015",
  "USGS:07103980:00011:00014",
  "USGS:07047942:00011:00002",
  "USGS:07047942:00011:00003",
  "USGS:07047950:00011:00001",
  "USGS:07047950:00011:00002",
  "USGS:07048480:00011:00002",
  "USGS:07048480:00011:00003",
  "USGS:07048480:00011:00001",
  "USGS:08405200:00011:00014",
  "USGS:08405200:00011:00001",
  "USGS:08405200:00011:00002",
  "USGS:08405200:00011:00015",
  "USGS:08405450:00011:00002",
  "USGS:08405450:00011:00001",
  "USGS:08405500:00011:00001",
  "USGS:08405500:00011:00002",
  "USGS:08406000:00011:00002",
  "USGS:08406000:00011:00001",
  "USGS:08406500:00011:00015",
  "USGS:08406500:00011:00002",
  "USGS:08406500:00011:00004",
  "USGS:08406500:00011:00016",
  "USGS:08407000:00011:00002",
  "USGS:08407000:00011:00004",
  "USGS:08407500:00011:00016",
  "USGS:08407500:00011:00001",
  "USGS:08407500:00011:00002",
  "USGS:08407500:00011:00017",
  "USGS:08408500:00011:00001",
  "USGS:08408500:00011:00002",
  "USGS:08477110:00011:00001",
  "USGS:08477110:00011:00002",
  "USGS:08481500:00011:00001",
  "USGS:08481500:00011:00002",
  "USGS:09355500:00011:00006",
  "USGS:09355500:00011:00007",
  "USGS:09355500:00011:00008",
  "USGS:09364010:00011:00002",
  "USGS:09364010:00011:00001",
  "USGS:09364500:00011:00002",
  "USGS:09364500:00011:00006",
  "USGS:09365000:00011:00016",
  "USGS:09365000:00011:00005",
  "USGS:09365000:00011:00006",
  "USGS:09367000:00011:00002",
  "USGS:09367000:00011:00001",
  "USGS:09367500:00011:00001",
  "USGS:09367500:00011:00002",
  "USGS:09367580:00011:00001",
  "USGS:09367580:00011:00002",
  "USGS:09367580:00011:00004",
  "USGS:09368000:00011:00008",
  "USGS:09368000:00011:00012",
  "USGS:09386900:00011:00001",
  "USGS:09386900:00011:00002",
  "USGS:09386950:00011:00001",
  "USGS:09386950:00011:00002",
  "USGS:09430500:00011:00005",
  "USGS:09430500:00011:00006",
  "USGS:09430600:00011:00001",
  "USGS:09430600:00011:00002",
  "USGS:09431500:00011:00005",
  "USGS:09431500:00011:00006",
  "USGS:09432000:00011:00001",
  "USGS:09432000:00011:00002",
  "USGS:09442680:00011:00001",
  "USGS:09442680:00011:00002",
  "USGS:09442980:00011:00005",
  "USGS:09442980:00011:00001",
  "USGS:09442980:00011:00003",
  "USGS:09443800:00011:00006",
  "USGS:09443800:00011:00001",
  "USGS:09443800:00011:00002",
  "USGS:09444000:00011:00005",
  "USGS:09444000:00011:00006",
  "USGS:321740106481001:00011:00001",
  "USGS:321740106481003:00011:00001",
  "USGS:321740106481004:00011:00001",
  "USGS:321745106492101:00011:00001",
  "USGS:321745106492102:00011:00001",
  "USGS:321745106492103:00011:00001",
  "USGS:321745106492106:00011:00001",
  "USGS:322323106314701:00011:00001",
  "USGS:323733107011002:00011:00003",
  "USGS:323733107011002:00011:00004",
  "USGS:323733107011002:00011:00006",
  "USGS:323733107011002:00011:00005",
  "USGS:323733107011002:00011:00001",
  "USGS:324007107095501:00011:00003",
  "USGS:324007107095501:00011:00004",
  "USGS:324007107095501:00011:00006",
  "USGS:324007107095501:00011:00005",
  "USGS:324007107095501:00011:00001",
  "USGS:324955107180902:00011:00003",
  "USGS:324955107180902:00011:00004",
  "USGS:324955107180902:00011:00006",
  "USGS:324955107180902:00011:00005",
  "USGS:324955107180902:00011:00001",
  "USGS:331421108484500:00011:00001",
  "USGS:331617108353900:00011:00001",
  "USGS:331950108383800:00011:00001",
  "USGS:332538105440401:00011:00001",
  "USGS:332538105440401:00011:00003",
  "USGS:332659108400700:00011:00001",
  "USGS:332748105481601:00011:00001",
  "USGS:332748105481601:00011:00003",
  "USGS:332940105470501:00011:00001",
  "USGS:332940105470501:00011:00003",
  "USGS:09022000:00011:00003",
  "USGS:09022000:00011:00005",
  "USGS:09024000:00011:00003",
  "USGS:09024000:00011:00002",
  "USGS:09025000:00011:00003",
  "USGS:09025000:00011:00014",
  "USGS:09025300:00011:00002",
  "USGS:09025300:00011:00001",
  "USGS:09026500:00011:00002",
  "USGS:09026500:00011:00004",
  "USGS:09027100:00011:00013",
  "USGS:09027100:00011:00002",
  "USGS:0204382800:00011:00017",
  "USGS:02053200:00011:00001",
  "USGS:02053200:00011:00002",
  "USGS:02053500:00011:00001",
  "USGS:02053500:00011:00002",
  "USGS:02068500:00011:00001",
  "USGS:02068500:00011:00002",
  "USGS:02069000:00011:00006",
  "USGS:02069000:00011:00001",
  "USGS:02069000:00011:00002",
  "USGS:02070500:00011:00002",
  "USGS:02070500:00011:00003",
  "USGS:02071000:00011:00002",
  "USGS:02071000:00011:00003",
  "USGS:02074000:00011:00002",
  "USGS:02074000:00011:00003",
  "USGS:02077200:00011:00001",
  "USGS:02077200:00011:00002",
  "USGS:02077200:00011:00003",
  "USGS:02077280:00011:00002",
  "USGS:02077280:00011:00012",
  "USGS:0207730290:00011:00001",
  "USGS:02077303:00011:00001",
  "USGS:02077303:00011:00002",
  "USGS:02077303:00011:00003",
  "USGS:02077670:00011:00001",
  "USGS:02077670:00011:00002",
  "USGS:02080500:00011:00004",
  "USGS:02080500:00011:00005",
  "USGS:0208062765:00011:00002",
  "USGS:0208062765:00011:00001",
  "USGS:0208062765:00011:00003",
  "USGS:0208062765:00011:00006",
  "USGS:0208062765:00011:00005",
  "USGS:0208062765:00011:00008",
  "USGS:02081000:00011:00006",
  "USGS:02081022:00011:00004",
  "USGS:02081022:00011:00003",
  "USGS:02081022:00011:00005",
  "USGS:02081022:00011:00008",
  "USGS:02081022:00011:00007",
  "USGS:02081022:00011:00010",
  "USGS:02081028:00011:00001",
  "USGS:340800117235903:00011:00001",
  "USGS:340800117235904:00011:00001",
  "USGS:340804117221601:00011:00001",
  "USGS:340804117221602:00011:00001",
  "USGS:340804117221603:00011:00001",
  "USGS:340804117221604:00011:00001",
  "USGS:341509117312601:00011:00001",
  "USGS:341512117102201:00011:00001",
  "USGS:341545117124001:00011:00001",
  "USGS:341602117110401:00011:00001",
  "USGS:342630119442301:00011:00003",
  "USGS:342630119442301:00011:00001",
  "USGS:343120118533301:00011:00001",
  "USGS:364200119420001:00011:00001",
  "USGS:364200119420001:00011:00002",
  "USGS:364200119420001:00011:00006",
  "USGS:364200119420001:00011:00005",
  "USGS:364200119420001:00011:00004",
  "USGS:364200119420001:00011:00003",
  "USGS:364200119420001:00011:00007",
  "USGS:373015122071000:00011:00010",
  "USGS:373015122071000:00011:00011",
  "USGS:373015122071000:00011:00020",
  "USGS:373015122071000:00011:00006",
  "USGS:373015122071000:00011:00007",
  "USGS:373015122071000:00011:00016",
  "USGS:373015122071000:00011:00017",
  "USGS:373015122071000:00011:00014",
  "USGS:373015122071000:00011:00015",
  "USGS:373015122071000:00011:00004",
  "USGS:373015122071000:00011:00005",
  "USGS:373025122065901:00011:00001",
  "USGS:373818118513301:00011:00002",
  "USGS:373818118513301:00011:00001",
  "USGS:373822118514401:00011:00006",
  "USGS:373822118514401:00011:00005",
  "USGS:373822118514401:00011:00004",
  "USGS:373822118514401:00011:00001",
  "USGS:373829118505801:00011:00003",
  "USGS:373829118505801:00011:00002",
  "USGS:373829118505801:00011:00001",
  "USGS:374811122235001:00011:00001",
  "USGS:374811122235001:00011:00002",
  "USGS:374811122235001:00011:00007",
  "USGS:374811122235001:00011:00006",
  "USGS:374811122235001:00011:00005",
  "USGS:374811122235001:00011:00003",
  "USGS:374938122251801:00011:00002",
  "USGS:374938122251801:00011:00001",
  "USGS:374938122251801:00011:00004",
  "USGS:374938122251801:00011:00005",
  "USGS:374938122251801:00011:00008",
  "USGS:375805121121101:00011:00001",
  "USGS:375805121121102:00011:00001",
  "USGS:375805121121103:00011:00001",
  "USGS:375805121121104:00011:00001",
  "USGS:385525122335501:00011:00001",
  "USGS:390500122321601:00011:00001",
  "USGS:390959120083601:00011:00013",
  "USGS:391056122420801:00011:00001",
  "USGS:391930120165301:00011:00005",
  "USGS:392541120015901:00011:00003",
  "USGS:392724120171001:00011:00002",
  "USGS:09143600:00011:00002",
  "USGS:09143600:00011:00001",
  "USGS:09144250:00011:00019",
  "USGS:09144250:00011:00001",
  "USGS:09144250:00011:00002",
  "USGS:09144250:00011:00021",
  "USGS:09146020:00011:00002",
  "USGS:09146020:00011:00001",
  "USGS:07076750:00011:00003",
  "USGS:07076750:00011:00006",
  "USGS:07076750:00011:00002",
  "USGS:07077000:00011:00002",
  "USGS:07077000:00011:00003",
  "USGS:07077380:00011:00016",
  "USGS:07077380:00011:00005",
  "USGS:07077380:00011:00004",
  "USGS:07077500:00011:00001",
  "USGS:07077555:00011:00011",
  "USGS:07077555:00011:00010",
  "USGS:07077652:00011:00002",
  "USGS:07077652:00011:00013",
  "USGS:07077652:00011:00001",
  "USGS:07077730:00011:00004",
  "USGS:07077730:00011:00003",
  "USGS:07077730:00011:00001",
  "USGS:07191160:00011:00003",
  "USGS:07191160:00011:00002",
  "USGS:07191160:00011:00001",
  "USGS:07191179:00011:00003",
  "USGS:07191179:00011:00002",
  "USGS:07191179:00011:00001",
  "USGS:07194800:00011:00001",
  "USGS:07194800:00011:00002",
  "USGS:07194809:00011:00002",
  "USGS:07194809:00011:00003",
  "USGS:07194809:00011:00001",
  "USGS:07194880:00011:00014",
  "USGS:07194880:00011:00012",
  "USGS:07194880:00011:00011",
  "USGS:07194880:00011:00001",
  "USGS:07194880:00011:00015",
  "USGS:07194880:00011:00016",
  "USGS:07194880:00011:00017",
  "USGS:07194906:00011:00005",
  "USGS:07194906:00011:00002",
  "USGS:07194906:00011:00001",
  "USGS:07194933:00011:00005",
  "USGS:07194933:00011:00003",
  "USGS:07194933:00011:00001",
  "USGS:07195000:00011:00002",
  "USGS:07195000:00011:00003",
  "USGS:07195400:00011:00004",
  "USGS:07195400:00011:00001",
  "USGS:07195400:00011:00002",
  "USGS:07195430:00011:00011",
  "USGS:07195430:00011:00001",
  "USGS:07195800:00011:00003",
  "USGS:07195800:00011:00004",
  "USGS:07196900:00011:00016",
  "USGS:07196900:00011:00005",
  "USGS:07196900:00011:00004",
  "USGS:07247000:00011:00015",
  "USGS:07247000:00011:00004",
  "USGS:07249400:00011:00002",
  "USGS:07249400:00011:00003",
  "USGS:07249455:00011:00015",
  "USGS:07249455:00011:00017",
  "USGS:07249455:00011:00001",
  "USGS:07250085:00011:00002",
  "USGS:07250085:00011:00012",
  "USGS:07250085:00011:00001",
  "USGS:07250550:00011:00001",
  "USGS:07250550:00011:00002",
  "USGS:07250550:00011:00003",
  "USGS:07250550:00011:00004",
  "USGS:07250550:00011:00005",
  "USGS:07250550:00011:00006",
  "USGS:07250550:00011:00007",
  "USGS:07250550:00011:00008",
  "USGS:07250550:00011:00009",
  "USGS:07250550:00011:00010",
  "USGS:07250550:00011:00011",
  "USGS:07250550:00011:00012",
  "USGS:07250550:00011:00013",
  "USGS:07250550:00011:00014",
  "USGS:07250550:00011:00015",
  "USGS:07250550:00011:00016",
  "USGS:07250550:00011:00017",
  "USGS:07250550:00011:00018",
  "USGS:07250935:00011:00002",
  "USGS:07250935:00011:00004",
  "USGS:07250935:00011:00001",
  "USGS:07250965:00011:00002",
  "USGS:07250965:00011:00004",
  "USGS:07250965:00011:00001",
  "USGS:07250974:00011:00002",
  "USGS:07250974:00011:00013",
  "USGS:07250974:00011:00001",
  "USGS:07251500:00011:00003",
  "USGS:07251500:00011:00002",
  "USGS:07252000:00011:00004",
  "USGS:07252000:00011:00002",
  "USGS:07252000:00011:00003",
  "USGS:07256500:00011:00003",
  "USGS:07256500:00011:00002",
  "USGS:07257006:00011:00003",
  "USGS:07257006:00011:00002",
  "USGS:07257006:00011:00001",
  "USGS:07257200:00011:00004",
  "USGS:07257200:00011:00002",
  "USGS:07257450:00011:00002",
  "USGS:07257450:00011:00001",
  "USGS:07257460:00011:00001",
  "USGS:07257460:00011:00002",
  "USGS:07257473:00011:00005",
  "USGS:07257473:00011:00001",
  "USGS:07257473:00011:00002",
  "USGS:07257480:00011:00002",
  "USGS:07257480:00011:00001",
  "USGS:07257500:00011:00004",
  "USGS:07257500:00011:00003",
  "USGS:07257500:00011:00005",
  "USGS:07257500:00011:00002",
  "USGS:07257500:00011:00006",
  "USGS:07257500:00011:00019",
  "USGS:07257500:00011:00017",
  "USGS:07257500:00011:00020",
  "USGS:07257500:00011:00018",
  "USGS:07257693:00011:00002",
  "USGS:07257693:00011:00014",
  "USGS:07257693:00011:00001",
  "USGS:07258000:00011:00007",
  "USGS:07258500:00011:00003",
  "USGS:07258500:00011:00005",
  "USGS:07258500:00011:00002",
  "USGS:07260000:00011:00003",
  "USGS:07260000:00011:00006",
  "USGS:07260000:00011:00002",
  "USGS:07260500:00011:00004",
  "USGS:07260500:00011:00002",
  "USGS:07260500:00011:00003",
  "USGS:07260640:00011:00003",
  "USGS:07260640:00011:00002",
  "USGS:09070000:00011:00001",
  "USGS:09070000:00011:00002",
  "USGS:09070500:00011:00001",
  "USGS:09070500:00011:00002",
  "USGS:09071750:00011:00004",
  "USGS:09071750:00011:00006",
  "USGS:09072550:00011:00001",
  "USGS:09072550:00011:00002",
  "USGS:09073005:00011:00001",
  "USGS:09073005:00011:00002",
  "USGS:09073300:00011:00001",
  "USGS:09073300:00011:00003",
  "USGS:09073400:00011:00001",
  "USGS:09073400:00011:00004",
  "USGS:09074000:00011:00004",
  "USGS:09074000:00011:00001",
  "USGS:09074500:00011:00002",
  "USGS:09074500:00011:00001",
  "USGS:06714360:00011:00001",
  "USGS:06714400:00011:00002",
  "USGS:06714400:00011:00001",
  "USGS:06714800:00011:00002",
  "USGS:06714800:00011:00001",
  "USGS:06715000:00011:00002",
  "USGS:06715000:00011:00004",
  "USGS:06716100:00011:00002",
  "USGS:06716100:00011:00004",
  "USGS:06716500:00011:00001",
  "USGS:06716500:00011:00002",
  "USGS:06718550:00011:00002",
  "USGS:06718550:00011:00001",
  "USGS:06719505:00011:00005",
  "USGS:06719505:00011:00003",
  "USGS:06719560:00011:00004",
  "USGS:06719560:00011:00003",
  "USGS:06719840:00011:00002",
  "USGS:06719840:00011:00001",
  "USGS:06720460:00011:00012",
  "USGS:06720460:00011:00002",
  "USGS:06720460:00011:00001",
  "USGS:06720820:00011:00002",
  "USGS:06720820:00011:00001",
  "USGS:06720990:00011:00002",
  "USGS:06720990:00011:00003",
  "USGS:06721000:00011:00001",
  "USGS:06721000:00011:00002",
  "USGS:06724970:00011:00002",
  "USGS:06724970:00011:00001",
  "USGS:06727500:00011:00001",
  "USGS:06727500:00011:00002",
  "USGS:06730160:00011:00002",
  "USGS:06730160:00011:00001",
  "USGS:06730160:00011:00003",
  "USGS:06730200:00011:00004",
  "USGS:06730200:00011:00003",
  "USGS:06730500:00011:00001",
  "USGS:06730500:00011:00002",
  "USGS:06730525:00011:00002",
  "USGS:06730525:00011:00001",
  "USGS:06741510:00011:00001",
  "USGS:06741510:00011:00002",
  "USGS:06746095:00011:00001",
  "USGS:06746095:00011:00003",
  "USGS:06746110:00011:00002",
  "USGS:06746110:00011:00001",
  "USGS:06751150:00011:00002",
  "USGS:06751150:00011:00001",
  "USGS:06751490:00011:00002",
  "USGS:06751490:00011:00006",
  "USGS:06752260:00011:00004",
  "USGS:06752260:00011:00002",
  "USGS:06752280:00011:00001",
  "USGS:06752280:00011:00002",
  "USGS:06759500:00011:00001",
  "USGS:06759500:00011:00002",
  "USGS:07079300:00011:00002",
  "USGS:07079300:00011:00008",
  "USGS:07081200:00011:00001",
  "USGS:07081200:00011:00006",
  "USGS:07083000:00011:00001",
  "USGS:07083000:00011:00005",
  "USGS:07083000:00011:00004",
  "USGS:07083200:00011:00001",
  "USGS:07083200:00011:00002",
  "USGS:07086000:00011:00012",
  "USGS:07086000:00011:00013",
  "USGS:07091200:00011:00003",
  "USGS:07091200:00011:00002",
  "USGS:07096000:00011:00003",
  "USGS:07096000:00011:00004",
  "USGS:07096250:00011:00004",
  "USGS:07096250:00011:00003",
  "USGS:07097000:00011:00017",
  "USGS:07097000:00011:00018",
  "USGS:07099050:00011:00002",
  "USGS:07099050:00011:00003",
  "USGS:07099060:00011:00013",
  "USGS:07099060:00011:00002",
  "USGS:07099060:00011:00003",
  "USGS:07099225:00011:00002",
  "USGS:07099225:00011:00001",
  "USGS:07099233:00011:00001",
  "USGS:07099233:00011:00003",
  "USGS:07099400:00011:00001",
  "USGS:07099400:00011:00003",
  "USGS:07363500:00011:00002",
  "USGS:07099969:00011:00004",
  "USGS:07099970:00011:00009",
  "USGS:07099970:00011:00021",
  "USGS:07099970:00011:00002",
  "USGS:07099970:00011:00008",
  "USGS:07099970:00011:00010",
  "USGS:07099973:00011:00002",
  "USGS:07099973:00011:00001",
  "USGS:07103700:00011:00001",
  "USGS:07103700:00011:00002",
  "USGS:07103700:00011:00003",
  "USGS:07103702:00011:00004",
  "USGS:07103702:00011:00002",
  "USGS:07103702:00011:00001",
  "USGS:07103703:00011:00014",
  "USGS:07103703:00011:00002",
  "USGS:07103703:00011:00001",
  "USGS:07103703:00011:00004",
  "USGS:09353800:00011:00002",
  "USGS:09353800:00011:00001",
  "USGS:09354500:00011:00001",
  "USGS:09354500:00011:00003",
  "USGS:09358000:00011:00013",
  "USGS:09358000:00011:00012",
  "USGS:09358550:00011:00004",
  "USGS:09358550:00011:00003",
  "USGS:09359010:00011:00004",
  "USGS:09359010:00011:00002",
  "USGS:09359020:00011:00008",
  "USGS:07360200:00011:00011",
  "USGS:07360200:00011:00001",
  "USGS:07361500:00011:00002",
  "USGS:07361500:00011:00003",
  "USGS:07362000:00011:00003",
  "USGS:07362000:00011:00006",
  "USGS:07362000:00011:00002",
  "USGS:07362100:00011:00002",
  "USGS:07362100:00011:00003",
  "USGS:07362500:00011:00002",
  "USGS:07362500:00011:00003",
  "USGS:07362579:00011:00002",
  "USGS:07362579:00011:00003",
  "USGS:07362579:00011:00004",
  "USGS:07362579:00011:00014",
  "USGS:07362579:00011:00001",
  "USGS:07362587:00011:00002",
  "USGS:07362587:00011:00001",
  "USGS:07362591:00011:00012",
  "USGS:07362591:00011:00013",
  "USGS:07362591:00011:00001",
  "USGS:07363000:00011:00005",
  "USGS:07363000:00011:00001",
  "USGS:07363000:00011:00004",
  "USGS:07363200:00011:00017",
  "USGS:07363200:00011:00001",
  "USGS:07363200:00011:00011",
  "USGS:07363400:00011:00004",
  "USGS:07363400:00011:00002",
  "USGS:07363400:00011:00001",
  "USGS:07363500:00011:00015",
  "USGS:07363500:00011:00003",
  "USGS:07364000:00011:00001",
  "USGS:07364078:00011:00002",
  "USGS:07364078:00011:00001",
  "USGS:07364122:00011:00006",
  "USGS:07364122:00011:00002",
  "USGS:07364122:00011:00005",
  "USGS:07364122:00011:00007",
  "USGS:07364130:00011:00006",
  "USGS:07364130:00011:00002",
  "USGS:07364130:00011:00003",
  "USGS:07364130:00011:00005",
  "USGS:07364130:00011:00007",
  "USGS:07364133:00011:00014",
  "USGS:07364133:00011:00002",
  "USGS:07364133:00011:00003",
  "USGS:07364150:00011:00003",
  "USGS:07364150:00011:00004",
  "USGS:07364185:00011:00016",
  "USGS:07364185:00011:00017",
  "USGS:07364185:00011:00001",
  "USGS:07367680:00011:00003",
  "USGS:07367680:00011:00001",
  "USGS:07369680:00011:00017",
  "USGS:07369680:00011:00003",
  "USGS:07369680:00011:00002",
  "USGS:07369680:00011:00001",
  "USGS:330624091552801:00011:00001",
  "USGS:331104092380201:00011:00001",
  "USGS:331256092483702:00011:00001",
  "USGS:331354092322401:00011:00001",
  "USGS:331438092411901:00011:00001",
  "USGS:331609093144902:00011:00001",
  "USGS:332205092433001:00011:00001",
  "USGS:335258091152301:00011:00001",
  "USGS:340747091214501:00011:00001",
  "USGS:340806091210701:00011:00001",
  "USGS:340859091211201:00011:00001",
  "USGS:341453091544101:00011:00001",
  "USGS:342649091251916:00011:00001",
  "USGS:343045093054901:00011:00001",
  "USGS:343048093030401:00011:00001",
  "USGS:343048093031301:00011:00001",
  "USGS:343049093031301:00011:00001",
  "USGS:343052093031301:00011:00001",
  "USGS:343054093031201:00011:00001",
  "USGS:343057093031301:00011:00001",
  "USGS:343108090462601:00011:00001",
  "USGS:343114930420001:00011:00001",
  "USGS:343204093005501:00011:00001",
  "USGS:343206093044101:00011:00001",
  "USGS:343255092593601:00011:00001",
  "USGS:01511000:00011:00003",
  "USGS:01511000:00011:00002",
  "USGS:01511000:00011:00001",
  "USGS:03086500:00011:00022",
  "USGS:03086500:00011:00003",
  "USGS:03090000:00011:00013",
  "USGS:03090500:00011:00015",
  "USGS:03090500:00011:00004",
  "USGS:06700000:00011:00013",
  "USGS:06700000:00011:00001",
  "USGS:06700000:00011:00002",
  "USGS:06701620:00011:00003",
  "USGS:06701620:00011:00002",
  "USGS:06701620:00011:00001",
  "USGS:06701700:00011:00013",
  "USGS:06701700:00011:00001",
  "USGS:06701900:00011:00002",
  "USGS:06701900:00011:00001",
  "USGS:06708600:00011:00002",
  "USGS:06708600:00011:00001",
  "USGS:06708800:00011:00002",
  "USGS:06708800:00011:00001",
  "USGS:06709000:00011:00003",
  "USGS:06709000:00011:00001",
  "USGS:06709000:00011:00002",
  "USGS:06709530:00011:00004",
  "USGS:06709530:00011:00001",
  "USGS:06709740:00011:00002",
  "USGS:06709740:00011:00001",
  "USGS:06709910:00011:00002",
  "USGS:06709910:00011:00001",
  "USGS:06710150:00011:00002",
  "USGS:06710150:00011:00001",
  "USGS:06710247:00011:00002",
  "USGS:06710247:00011:00001",
  "USGS:06710385:00011:00001",
  "USGS:06710385:00011:00004",
  "USGS:06710605:00011:00002",
  "USGS:06710605:00011:00005",
  "USGS:06711515:00011:00002",
  "USGS:06711515:00011:00001",
  "USGS:06711555:00011:00002",
  "USGS:06711555:00011:00001",
  "USGS:06711565:00011:00009",
  "USGS:06711565:00011:00002",
  "USGS:06711565:00011:00008",
  "USGS:06711565:00011:00010",
  "USGS:06711565:00011:00011",
  "USGS:06711565:00011:00012",
  "USGS:06711570:00011:00002",
  "USGS:06711570:00011:00003",
  "USGS:06711575:00011:00006",
  "USGS:06711575:00011:00004",
  "USGS:06711575:00011:00005",
  "USGS:06711618:00011:00002",
  "USGS:06711618:00011:00001",
  "USGS:06711770:00011:00002",
  "USGS:06711770:00011:00001",
  "USGS:06711780:00011:00002",
  "USGS:06711780:00011:00001",
  "USGS:06712000:00011:00007",
  "USGS:06712000:00011:00001",
  "USGS:06712000:00011:00005",
  "USGS:06713000:00011:00001",
  "USGS:06713000:00011:00004",
  "USGS:343312093013201:00011:00001",
  "USGS:343330092591101:00011:00001",
  "USGS:343350093005901:00011:00001",
  "USGS:343518092591701:00011:00001",
  "USGS:343726093481801:00011:00001",
  "USGS:344651091355102:00011:00001",
  "USGS:344653091382701:00011:00001",
  "USGS:345057091525601:00011:00003",
  "USGS:351354092232401:00011:00001",
  "USGS:352341090213101:00011:00001",
  "USGS:352644091110901:00011:00001",
  "USGS:352726090523101:00011:00002",
  "USGS:352828091114401:00011:00001",
  "USGS:353151091180301:00011:00001",
  "USGS:353219091163601:00011:00001",
  "USGS:353606090510701:00011:00001",
  "USGS:354048091035401:00011:00001",
  "USGS:354207091041901:00011:00001",
  "USGS:354252091042201:00011:00001",
  "USGS:354717091081701:00011:00001",
  "USGS:354916090512501:00011:00001",
  "USGS:355927092122401:00011:00001",
  "USGS:07148400:00011:00016",
  "USGS:07148400:00011:00006",
  "USGS:07148400:00011:00005",
  "USGS:07149520:00011:00001",
  "USGS:07149520:00011:00004",
  "USGS:07151000:00011:00014",
  "USGS:07151000:00011:00013",
  "USGS:07151000:00011:00012",
  "USGS:07260672:00011:00003",
  "USGS:07260672:00011:00001",
  "USGS:07260673:00011:00013",
  "USGS:07260673:00011:00002",
  "USGS:07260678:00011:00002",
  "USGS:07260678:00011:00005",
  "USGS:07260678:00011:00001",
  "USGS:07260800:00011:00003",
  "USGS:07260800:00011:00002",
  "USGS:07260990:00011:00005",
  "USGS:07260990:00011:00002",
  "USGS:07260990:00011:00007",
  "USGS:07260990:00011:00001",
  "USGS:07261000:00011:00013",
  "USGS:07261000:00011:00001",
  "USGS:07261000:00011:00002",
  "USGS:07261090:00011:00004",
  "USGS:07261090:00011:00005",
  "USGS:07261090:00011:00003",
  "USGS:07261090:00011:00002",
  "USGS:07261090:00011:00001",
  "USGS:07261090:00011:00019",
  "USGS:07261090:00011:00016",
  "USGS:07261090:00011:00017",
  "USGS:07261090:00011:00018",
  "USGS:07261090:00011:00020",
  "USGS:07261200:00011:00001",
  "USGS:07261250:00011:00019",
  "USGS:07261250:00011:00021",
  "USGS:07261250:00011:00022",
  "USGS:07261250:00011:00017",
  "USGS:07261500:00011:00004",
  "USGS:07261500:00011:00002",
  "USGS:07261500:00011:00003",
  "USGS:07263000:00011:00003",
  "USGS:07263000:00011:00002",
  "USGS:07263012:00011:00003",
  "USGS:07263012:00011:00012",
  "USGS:07263012:00011:00002",
  "USGS:07263295:00011:00014",
  "USGS:07263295:00011:00002",
  "USGS:07263295:00011:00001",
  "USGS:07263296:00011:00013",
  "USGS:07263296:00011:00002",
  "USGS:07263296:00011:00001",
  "USGS:07263296:00011:00015",
  "USGS:07263296:00011:00014",
  "USGS:07263296:00011:00017",
  "USGS:07263296:00011:00018",
  "USGS:07263296:00011:00020",
  "USGS:072632962:00011:00003",
  "USGS:072632962:00011:00002",
  "USGS:072632962:00011:00001",
  "USGS:072632966:00011:00023",
  "USGS:072632966:00011:00002",
  "USGS:072632966:00011:00004",
  "USGS:072632966:00011:00009",
  "USGS:072632966:00011:00019",
  "USGS:072632966:00011:00001",
  "USGS:072632966:00011:00017",
  "USGS:072632966:00011:00020",
  "USGS:072632966:00011:00021",
  "USGS:072632966:00011:00022",
  "USGS:072632968:00011:00003",
  "USGS:072632968:00011:00002",
  "USGS:072632968:00011:00005",
  "USGS:072632968:00011:00001",
  "USGS:072632971:00011:00002",
  "USGS:072632971:00011:00001",
  "USGS:072632982:00011:00002",
  "USGS:072632982:00011:00001",
  "USGS:072632995:00011:00010",
  "USGS:072632995:00011:00011",
  "USGS:072632995:00011:00012",
  "USGS:072632995:00011:00013",
  "USGS:072632995:00011:00014",
  "USGS:072632995:00011:00015",
  "USGS:072632995:00011:00016",
  "USGS:072632995:00011:00018",
  "USGS:072632995:00011:00048",
  "USGS:072632995:00011:00049",
  "USGS:072632995:00011:00050",
  "USGS:072632995:00011:00051",
  "USGS:072632995:00011:00025",
  "USGS:072632995:00011:00021",
  "USGS:072632995:00011:00020",
  "USGS:072632995:00011:00024",
  "USGS:072632995:00011:00001",
  "USGS:072632995:00011:00002",
  "USGS:072632995:00011:00003",
  "USGS:072632995:00011:00004",
  "USGS:072632995:00011:00005",
  "USGS:072632995:00011:00006",
  "USGS:072632995:00011:00007",
  "USGS:072632995:00011:00009",
  "USGS:072632995:00011:00047",
  "USGS:072632995:00011:00052",
  "USGS:072632995:00011:00053",
  "USGS:072632995:00011:00054",
  "USGS:072632995:00011:00023",
  "USGS:072632995:00011:00045",
  "USGS:072632995:00011:00019",
  "USGS:072632995:00011:00022",
  "USGS:07263300:00011:00013",
  "USGS:07263300:00011:00012",
  "USGS:07263300:00011:00001",
  "USGS:07263450:00011:00004",
  "USGS:07263450:00011:00002",
  "USGS:07263450:00011:00003",
  "USGS:07263450:00011:00022",
  "USGS:07263450:00011:00023",
  "USGS:07263450:00011:00024",
  "USGS:07263450:00011:00025",
  "USGS:07263450:00011:00026",
  "USGS:07263450:00011:00027",
  "USGS:07263450:00011:00028",
  "USGS:07263450:00011:00029",
  "USGS:07263450:00011:00030",
  "USGS:07263450:00011:00031",
  "USGS:07263450:00011:00032",
  "USGS:07263450:00011:00033",
  "USGS:07263450:00011:00034",
  "USGS:07263450:00011:00035",
  "USGS:07263500:00011:00002",
  "USGS:07263555:00011:00005",
  "USGS:07263555:00011:00004",
  "USGS:07263555:00011:00002",
  "USGS:07263555:00011:00001",
  "USGS:07263580:00011:00002",
  "USGS:07263580:00011:00001",
  "USGS:07263605:00011:00005",
  "USGS:07263605:00011:00003",
  "USGS:07263605:00011:00002",
  "USGS:07263605:00011:00001",
  "USGS:07263650:00011:00001",
  "USGS:07264000:00011:00002",
  "USGS:07264000:00011:00003",
  "USGS:07265280:00011:00001",
  "USGS:07337000:00011:00005",
  "USGS:07337000:00011:00004",
  "USGS:07337000:00011:00002",
  "USGS:07337000:00011:00003",
  "USGS:07339500:00011:00003",
  "USGS:07339500:00011:00002",
  "USGS:07340000:00011:00004",
  "USGS:07340000:00011:00002",
  "USGS:07340000:00011:00003",
  "USGS:07340300:00011:00014",
  "USGS:07340300:00011:00002",
  "USGS:07340300:00011:00004",
  "USGS:07340500:00011:00004",
  "USGS:07340500:00011:00002",
  "USGS:07341000:00011:00003",
  "USGS:07341000:00011:00002",
  "USGS:07341200:00011:00004",
  "USGS:07341200:00011:00002",
  "USGS:07341200:00011:00003",
  "USGS:07344370:00011:00011",
  "USGS:07344370:00011:00001",
  "USGS:07344370:00011:00013",
  "USGS:07355860:00011:00001",
  "USGS:07355870:00011:00002",
  "USGS:07355880:00011:00005",
  "USGS:07355880:00011:00004",
  "USGS:07355880:00011:00002",
  "USGS:07355880:00011:00006",
  "USGS:07355880:00011:00007",
  "USGS:07356000:00011:00002",
  "USGS:07356000:00011:00003",
  "USGS:07358250:00011:00001",
  "USGS:07358250:00011:00002",
  "USGS:07358250:00011:00003",
  "USGS:07358253:00011:00002",
  "USGS:07358253:00011:00003",
  "USGS:07358253:00011:00001",
  "USGS:07358257:00011:00003",
  "USGS:07358257:00011:00002",
  "USGS:07358257:00011:00001",
  "USGS:07358280:00011:00001",
  "USGS:07358280:00011:00029",
  "USGS:07358280:00011:00025",
  "USGS:07358280:00011:00024",
  "USGS:07358280:00011:00028",
  "USGS:07358280:00011:00003",
  "USGS:07358280:00011:00002",
  "USGS:07358280:00011:00004",
  "USGS:07358280:00011:00006",
  "USGS:07358280:00011:00027",
  "USGS:07358280:00011:00030",
  "USGS:07358280:00011:00026",
  "USGS:07358284:00011:00013",
  "USGS:07358284:00011:00003",
  "USGS:07358284:00011:00002",
  "USGS:405051083391201:00011:00004",
  "USGS:405051083391201:00011:00002",
  "USGS:405051083391201:00011:00001",
  "USGS:405051083391201:00011:00009",
  "USGS:405051083391201:00011:00005",
  "USGS:405209082393200:00011:00001",
  "USGS:03127000:00011:00003",
  "USGS:03127500:00011:00003",
  "USGS:03128500:00011:00003",
  "USGS:03129000:00011:00003",
  "USGS:03129000:00011:00001",
  "USGS:03129197:00011:00011",
  "USGS:03129197:00011:00001",
  "USGS:03130000:00011:00003",
  "USGS:03131500:00011:00007",
  "USGS:03133500:00011:00003",
  "USGS:03135000:00011:00003",
  "USGS:03136500:00011:00017",
  "USGS:03158200:00011:00003",
  "USGS:09075400:00011:00012",
  "USGS:09075400:00011:00002",
  "USGS:09075400:00011:00001",
  "USGS:09078475:00011:00002",
  "USGS:09078475:00011:00001",
  "USGS:09079450:00011:00002",
  "USGS:09079450:00011:00001",
  "USGS:09080400:00011:00014",
  "USGS:09080400:00011:00002",
  "USGS:09081000:00011:00002",
  "USGS:09081000:00011:00001",
  "USGS:09081600:00011:00001",
  "USGS:09081600:00011:00002",
  "USGS:09085000:00011:00004",
  "USGS:09085000:00011:00001",
  "USGS:09085000:00011:00002",
  "USGS:09085100:00011:00001",
  "USGS:09085100:00011:00004",
  "USGS:09085150:00011:00001",
  "USGS:09085150:00011:00002",
  "USGS:09091900:00011:00003",
  "USGS:09091900:00011:00002",
  "USGS:09091900:00011:00001",
  "USGS:09095500:00011:00004",
  "USGS:09095500:00011:00001",
  "USGS:09095500:00011:00002",
  "USGS:09095500:00011:00006",
  "USGS:09096100:00011:00003",
  "USGS:09096100:00011:00002",
  "USGS:09096100:00011:00004",
  "USGS:09096100:00011:00005",
  "USGS:09096100:00011:00001",
  "USGS:09096570:00011:00003",
  "USGS:09096570:00011:00013",
  "USGS:09096600:00011:00013",
  "USGS:09096600:00011:00001",
  "USGS:09105000:00011:00016",
  "USGS:09105000:00011:00006",
  "USGS:09105000:00011:00005",
  "USGS:09105000:00011:00018",
  "USGS:09106150:00011:00015",
  "USGS:09106150:00011:00014",
  "USGS:09107000:00011:00013",
  "USGS:09107000:00011:00003",
  "USGS:09109000:00011:00004",
  "USGS:09109000:00011:00006",
  "USGS:09109000:00011:00005",
  "USGS:09110000:00011:00001",
  "USGS:09110000:00011:00002",
  "USGS:09111250:00011:00002",
  "USGS:09111250:00011:00001",
  "USGS:09112200:00011:00001",
  "USGS:09112200:00011:00002",
  "USGS:09112500:00011:00001",
  "USGS:09112500:00011:00004",
  "USGS:09113980:00011:00001",
  "USGS:09113980:00011:00002",
  "USGS:09114500:00011:00001",
  "USGS:09114500:00011:00002",
  "USGS:09115500:00011:00001",
  "USGS:09115500:00011:00004",
  "USGS:09118450:00011:00001",
  "USGS:09118450:00011:00003",
  "USGS:09119000:00011:00004",
  "USGS:09119000:00011:00001",
  "USGS:09119000:00011:00003",
  "USGS:09123450:00011:00002",
  "USGS:09123450:00011:00001",
  "USGS:09124500:00011:00001",
  "USGS:09124500:00011:00003",
  "USGS:09125800:00011:00002",
  "USGS:09125800:00011:00001",
  "USGS:09126000:00011:00001",
  "USGS:09126000:00011:00002",
  "USGS:09127000:00011:00001",
  "USGS:09127000:00011:00002",
  "USGS:09128000:00011:00004",
  "USGS:09128000:00011:00003",
  "USGS:09129550:00011:00002",
  "USGS:09129550:00011:00001",
  "USGS:09129600:00011:00001",
  "USGS:09129600:00011:00002",
  "USGS:09129600:00011:00003",
  "USGS:09131495:00011:00004",
  "USGS:09131495:00011:00003",
  "USGS:09131495:00011:00002",
  "USGS:09131495:00011:00001",
  "USGS:09132500:00011:00001",
  "USGS:09132500:00011:00002",
  "USGS:09134100:00011:00002",
  "USGS:09134100:00011:00001",
  "USGS:09136100:00011:00003",
  "USGS:09136100:00011:00002",
  "USGS:09136100:00011:00001",
  "USGS:09136100:00011:00004",
  "USGS:09143000:00011:00001",
  "USGS:09143000:00011:00002",
  "USGS:09143500:00011:00001",
  "USGS:09143500:00011:00002",
  "USGS:03205470:00011:00002",
  "USGS:03205470:00011:00001",
  "USGS:03217200:00011:00001",
  "USGS:03217500:00011:00013",
  "USGS:03217500:00011:00002",
  "USGS:03217500:00011:00001",
  "USGS:03219500:00011:00001",
  "USGS:03219500:00011:00007",
  "USGS:03219500:00011:00006",
  "USGS:03219500:00011:00019",
  "USGS:03219500:00011:00020",
  "USGS:03219500:00011:00022",
  "USGS:03220000:00011:00005",
  "USGS:03220000:00011:00004",
  "USGS:03220500:00011:00003",
  "USGS:03220510:00011:00001",
  "USGS:03220510:00011:00002",
  "USGS:03220510:00011:00003",
  "USGS:03220510:00011:00004",
  "USGS:03221000:00011:00004",
  "USGS:03221000:00011:00003",
  "USGS:07103980:00011:00002",
  "USGS:07103980:00011:00004",
  "USGS:07103990:00011:00001",
  "USGS:07103990:00011:00012",
  "USGS:07103990:00011:00014",
  "USGS:07103990:00011:00015",
  "USGS:07104000:00011:00004",
  "USGS:07104000:00011:00003",
  "USGS:07104905:00011:00004",
  "USGS:07104905:00011:00003",
  "USGS:07104905:00011:00002",
  "USGS:07104905:00011:00015",
  "USGS:07104905:00011:00016",
  "USGS:07105000:00011:00015",
  "USGS:07105000:00011:00002",
  "USGS:07105000:00011:00005",
  "USGS:07105490:00011:00005",
  "USGS:07105490:00011:00002",
  "USGS:07105490:00011:00001",
  "USGS:07105500:00011:00004",
  "USGS:07105500:00011:00003",
  "USGS:07105500:00011:00018",
  "USGS:07105500:00011:00019",
  "USGS:07105530:00011:00004",
  "USGS:07105530:00011:00003",
  "USGS:07105600:00011:00015",
  "USGS:07105600:00011:00002",
  "USGS:07105600:00011:00001",
  "USGS:07105800:00011:00028",
  "USGS:07105800:00011:00004",
  "USGS:07105800:00011:00003",
  "USGS:07105800:00011:00026",
  "USGS:07105800:00011:00027",
  "USGS:07105900:00011:00001",
  "USGS:07105900:00011:00003",
  "USGS:07105940:00011:00001",
  "USGS:07105940:00011:00002",
  "USGS:07105940:00011:00013",
  "USGS:07105940:00011:00014",
  "USGS:07105945:00011:00001",
  "USGS:07105945:00011:00005",
  "USGS:07106000:00011:00018",
  "USGS:07106000:00011:00004",
  "USGS:07106000:00011:00003",
  "USGS:07106000:00011:00019",
  "USGS:07106000:00011:00021",
  "USGS:07106000:00011:00020",
  "USGS:07106300:00011:00001",
  "USGS:07106300:00011:00002",
  "USGS:07106500:00011:00019",
  "USGS:07106500:00011:00006",
  "USGS:07106500:00011:00002",
  "USGS:07106500:00011:00005",
  "USGS:07106500:00011:00020",
  "USGS:07106500:00011:00004",
  "USGS:07106500:00011:00021",
  "USGS:07108900:00011:00004",
  "USGS:07108900:00011:00003",
  "USGS:07109500:00011:00007",
  "USGS:07109500:00011:00001",
  "USGS:07109500:00011:00002",
  "USGS:07109500:00011:00008",
  "USGS:07109500:00011:00023",
  "USGS:07109500:00011:00022",
  "USGS:07116500:00011:00001",
  "USGS:07116500:00011:00003",
  "USGS:07119500:00011:00002",
  "USGS:07119500:00011:00005",
  "USGS:07119700:00011:00003",
  "USGS:07119700:00011:00004",
  "USGS:07120500:00011:00016",
  "USGS:07120500:00011:00017",
  "USGS:07121500:00011:00004",
  "USGS:07121500:00011:00003",
  "USGS:07124000:00011:00015",
  "USGS:07124000:00011:00001",
  "USGS:07124000:00011:00002",
  "USGS:07124000:00011:00016",
  "USGS:07124200:00011:00008",
  "USGS:07124200:00011:00007",
  "USGS:07124400:00011:00004",
  "USGS:07124400:00011:00003",
  "USGS:07124410:00011:00006",
  "USGS:07124410:00011:00005",
  "USGS:07126200:00011:00017",
  "USGS:07126200:00011:00002",
  "USGS:07126200:00011:00005",
  "USGS:07126300:00011:00001",
  "USGS:07126300:00011:00002",
  "USGS:07126480:00011:00009",
  "USGS:07126480:00011:00002",
  "USGS:07126480:00011:00007",
  "USGS:07126480:00011:00004",
  "USGS:07126480:00011:00005",
  "USGS:07126485:00011:00009",
  "USGS:07126485:00011:00008",
  "USGS:07128500:00011:00001",
  "USGS:07128500:00011:00002",
  "USGS:07130000:00011:00012",
  "USGS:07130000:00011:00001",
  "USGS:07130500:00011:00015",
  "USGS:07130500:00011:00001",
  "USGS:07130500:00011:00002",
  "USGS:07130500:00011:00016",
  "USGS:07133000:00011:00001",
  "USGS:07133000:00011:00006",
  "USGS:07134100:00011:00014",
  "USGS:07134100:00011:00001",
  "USGS:07134100:00011:00002",
  "USGS:07134180:00011:00004",
  "USGS:07134180:00011:00003",
  "USGS:07134990:00011:00002",
  "USGS:07134990:00011:00001",
  "USGS:08227000:00011:00004",
  "USGS:08261000:00011:00001",
  "USGS:08261000:00011:00002",
  "USGS:09010500:00011:00001",
  "USGS:09010500:00011:00005",
  "USGS:09027100:00011:00001",
  "USGS:09014050:00011:00008",
  "USGS:09014050:00011:00002",
  "USGS:09014050:00011:00006",
  "USGS:09014050:00011:00001",
  "USGS:09014050:00011:00010",
  "USGS:09014050:00011:00013",
  "USGS:09014050:00011:00012",
  "USGS:09014050:00011:00014",
  "USGS:09014050:00011:00011",
  "USGS:09015000:00011:00002",
  "USGS:09019500:00011:00001",
  "USGS:09019500:00011:00003",
  "USGS:404440074211301:00011:00002",
  "USGS:03245500:00011:00007",
  "USGS:03245500:00011:00006",
  "USGS:03246500:00011:00001",
  "USGS:03246500:00011:00002",
  "USGS:03247040:00011:00001",
  "USGS:03247041:00011:00005",
  "USGS:03247041:00011:00002",
  "USGS:03247500:00011:00003",
  "USGS:03247500:00011:00001",
  "USGS:03255000:00011:00001",
  "USGS:03255300:00011:00002",
  "USGS:03255300:00011:00001",
  "USGS:03255349:00011:00001",
  "USGS:03255390:00011:00002",
  "USGS:03255390:00011:00001",
  "USGS:03255420:00011:00002",
  "USGS:09032000:00011:00015",
  "USGS:09032000:00011:00001",
  "USGS:09032000:00011:00005",
  "USGS:09032100:00011:00001",
  "USGS:09032100:00011:00003",
  "USGS:09033100:00011:00013",
  "USGS:09033100:00011:00002",
  "USGS:09033100:00011:00003",
  "USGS:09033300:00011:00013",
  "USGS:09033300:00011:00002",
  "USGS:09033300:00011:00003",
  "USGS:09034250:00011:00001",
  "USGS:09034250:00011:00004",
  "USGS:09034900:00011:00001",
  "USGS:09034900:00011:00004",
  "USGS:09035500:00011:00001",
  "USGS:09035500:00011:00004",
  "USGS:09035700:00011:00001",
  "USGS:09035700:00011:00004",
  "USGS:09035900:00011:00001",
  "USGS:09035900:00011:00003",
  "USGS:09036000:00011:00001",
  "USGS:09036000:00011:00003",
  "USGS:09037500:00011:00002",
  "USGS:09037500:00011:00006",
  "USGS:09038500:00011:00002",
  "USGS:09038500:00011:00005",
  "USGS:09041090:00011:00014",
  "USGS:09041090:00011:00002",
  "USGS:09066200:00011:00001",
  "USGS:09041090:00011:00001",
  "USGS:09041090:00011:00015",
  "USGS:09041395:00011:00002",
  "USGS:09041395:00011:00001",
  "USGS:09041400:00011:00003",
  "USGS:09041400:00011:00002",
  "USGS:09041400:00011:00001",
  "USGS:09041400:00011:00004",
  "USGS:09041400:00011:00005",
  "USGS:09041900:00011:00001",
  "USGS:09041900:00011:00004",
  "USGS:09044300:00011:00001",
  "USGS:09044300:00011:00004",
  "USGS:09044800:00011:00001",
  "USGS:09044800:00011:00004",
  "USGS:09046490:00011:00001",
  "USGS:09046490:00011:00004",
  "USGS:09046600:00011:00001",
  "USGS:09046600:00011:00003",
  "USGS:09047500:00011:00001",
  "USGS:09047500:00011:00002",
  "USGS:09047700:00011:00001",
  "USGS:09047700:00011:00005",
  "USGS:09050100:00011:00001",
  "USGS:09050100:00011:00002",
  "USGS:09050700:00011:00004",
  "USGS:09050700:00011:00003",
  "USGS:09051050:00011:00002",
  "USGS:09051050:00011:00005",
  "USGS:09056500:00011:00006",
  "USGS:09056500:00011:00004",
  "USGS:09056500:00011:00005",
  "USGS:09056500:00011:00007",
  "USGS:09056500:00011:00002",
  "USGS:09056500:00011:00001",
  "USGS:09056500:00011:00017",
  "USGS:09057500:00011:00005",
  "USGS:09057500:00011:00002",
  "USGS:09058000:00011:00016",
  "USGS:09058000:00011:00005",
  "USGS:09058000:00011:00002",
  "USGS:09058500:00011:00001",
  "USGS:09058500:00011:00004",
  "USGS:09059500:00011:00004",
  "USGS:09059500:00011:00003",
  "USGS:09061600:00011:00002",
  "USGS:09061600:00011:00001",
  "USGS:09063000:00011:00007",
  "USGS:09063000:00011:00006",
  "USGS:09064000:00011:00001",
  "USGS:09064000:00011:00003",
  "USGS:09064600:00011:00002",
  "USGS:09064600:00011:00003",
  "USGS:09065100:00011:00001",
  "USGS:09065100:00011:00003",
  "USGS:09065500:00011:00001",
  "USGS:09065500:00011:00004",
  "USGS:09066000:00011:00001",
  "USGS:09066000:00011:00003",
  "USGS:09066200:00011:00004",
  "USGS:09066300:00011:00001",
  "USGS:09066300:00011:00003",
  "USGS:09066325:00011:00002",
  "USGS:09066325:00011:00001",
  "USGS:09066510:00011:00013",
  "USGS:09066510:00011:00002",
  "USGS:09066510:00011:00001",
  "USGS:09067000:00011:00001",
  "USGS:09067000:00011:00005",
  "USGS:09067020:00011:00002",
  "USGS:09067020:00011:00001",
  "USGS:09067200:00011:00001",
  "USGS:09067200:00011:00004",
  "USGS:04185440:00011:00002",
  "USGS:04185440:00011:00001",
  "USGS:04186500:00011:00002",
  "USGS:04186500:00011:00007",
  "USGS:04187100:00011:00002",
  "USGS:04187100:00011:00001",
  "USGS:04188100:00011:00002",
  "USGS:04188100:00011:00003",
  "USGS:04188337:00011:00003",
  "USGS:04188337:00011:00002",
  "USGS:04188337:00011:00001",
  "USGS:04188400:00011:00003",
  "USGS:04188400:00011:00002",
  "USGS:04188400:00011:00001",
  "USGS:04188433:00011:00003",
  "USGS:04188433:00011:00002",
  "USGS:09359020:00011:00007",
  "USGS:09359080:00011:00002",
  "USGS:09359080:00011:00001",
  "USGS:09359082:00011:00002",
  "USGS:09359082:00011:00001",
  "USGS:09359500:00011:00001",
  "USGS:09359500:00011:00002",
  "USGS:09361500:00011:00001",
  "USGS:09361500:00011:00002",
  "USGS:09362520:00011:00001",
  "USGS:09362520:00011:00002",
  "USGS:09362800:00011:00002",
  "USGS:09362800:00011:00001",
  "USGS:09363500:00011:00004",
  "USGS:09363500:00011:00005",
  "USGS:09370600:00011:00005",
  "USGS:09370600:00011:00004",
  "USGS:09371000:00011:00001",
  "USGS:09371000:00011:00005",
  "USGS:09371010:00011:00015",
  "USGS:09371010:00011:00001",
  "USGS:09371010:00011:00002",
  "USGS:09371492:00011:00003",
  "USGS:09371492:00011:00001",
  "USGS:09371492:00011:00002",
  "USGS:09371492:00011:00004",
  "USGS:09371520:00011:00003",
  "USGS:09371520:00011:00006",
  "USGS:09371520:00011:00005",
  "USGS:09371520:00011:00004",
  "USGS:09372000:00011:00001",
  "USGS:09372000:00011:00005",
  "USGS:351741080475045:00011:00004",
  "USGS:372319104073301:00011:00001",
  "USGS:372319104073301:00011:00005",
  "USGS:372319104073301:00011:00006",
  "USGS:372319104073301:00011:00013",
  "USGS:372319104073301:00011:00002",
  "USGS:372319104073301:00011:00003",
  "USGS:372319104073301:00011:00004",
  "USGS:372721103595601:00011:00001",
  "USGS:372721103595601:00011:00005",
  "USGS:372721103595601:00011:00011",
  "USGS:372721103595601:00011:00002",
  "USGS:372721103595601:00011:00003",
  "USGS:372721103595601:00011:00004",
  "USGS:373232103555201:00011:00001",
  "USGS:373232103555201:00011:00005",
  "USGS:373232103555201:00011:00011",
  "USGS:373232103555201:00011:00002",
  "USGS:373232103555201:00011:00003",
  "USGS:373232103555201:00011:00004",
  "USGS:373315103493101:00011:00001",
  "USGS:373315103493101:00011:00005",
  "USGS:373315103493101:00011:00011",
  "USGS:373315103493101:00011:00002",
  "USGS:373315103493101:00011:00003",
  "USGS:373315103493101:00011:00004",
  "USGS:373823103465601:00011:00001",
  "USGS:373823103465601:00011:00005",
  "USGS:373823103465601:00011:00011",
  "USGS:373823103465601:00011:00002",
  "USGS:373823103465601:00011:00003",
  "USGS:373823103465601:00011:00004",
  "USGS:374557105372401:00011:00002",
  "USGS:374557105372401:00011:00003",
  "USGS:374557105372401:00011:00004",
  "USGS:374557105372401:00011:00005",
  "USGS:374557105372401:00011:00001",
  "USGS:375546107412000:00011:00001",
  "USGS:375852107455200:00011:00001",
  "USGS:380251107513000:00011:00001",
  "USGS:380436107411500:00011:00001",
  "USGS:381312104321001:00011:00001",
  "USGS:381312104321001:00011:00002",
  "USGS:381312104321001:00011:00003",
  "USGS:382323104200701:00011:00011",
  "USGS:382323104200701:00011:00001",
  "USGS:382628104493700:00011:00002",
  "USGS:382628104493700:00011:00001",
  "USGS:382629104493000:00011:00002",
  "USGS:382629104493000:00011:00001",
  "USGS:383159104540701:00011:00001",
  "USGS:383159104540701:00011:00005",
  "USGS:383159104540701:00011:00011",
  "USGS:383159104540701:00011:00002",
  "USGS:383159104540701:00011:00003",
  "USGS:383159104540701:00011:00004",
  "USGS:383619104520401:00011:00002",
  "USGS:383619104520401:00011:00001",
  "USGS:383637104531301:00011:00002",
  "USGS:383637104531301:00011:00001",
  "USGS:383944104474201:00011:00002",
  "USGS:383944104474201:00011:00001",
  "USGS:383946107595301:00011:00002",
  "USGS:383946107595301:00011:00001",
  "USGS:384037104472001:00011:00002",
  "USGS:384037104472001:00011:00001",
  "USGS:384047104510301:00011:00002",
  "USGS:384047104510301:00011:00001",
  "USGS:384048104504901:00011:00002",
  "USGS:384048104504901:00011:00001",
  "USGS:384053104492001:00011:00001",
  "USGS:384053104492001:00011:00005",
  "USGS:384053104492001:00011:00011",
  "USGS:384053104492001:00011:00002",
  "USGS:384053104492001:00011:00003",
  "USGS:384053104492001:00011:00004",
  "USGS:384220104503701:00011:00002",
  "USGS:384220104503701:00011:00001",
  "USGS:384537104494701:00011:00002",
  "USGS:384908104453301:00011:00002",
  "USGS:384936107571901:00011:00001",
  "USGS:384936107571901:00011:00012",
  "USGS:384945107553401:00011:00001",
  "USGS:385010104422901:00011:00002",
  "USGS:385106106571000:00011:00002",
  "USGS:385106106571000:00011:00001",
  "USGS:04209000:00011:00007",
  "USGS:04209000:00011:00002",
  "USGS:04212100:00011:00020",
  "USGS:04212100:00011:00019",
  "USGS:04213000:00011:00017",
  "USGS:04213000:00011:00004",
  "USGS:04213000:00011:00003",
  "USGS:383638082103300:00011:00001",
  "USGS:390735084333300:00011:00003",
  "USGS:390735084333300:00011:00018",
  "USGS:390735084333300:00011:00017",
  "USGS:390735084333300:00011:00010",
  "USGS:390735084333300:00011:00011",
  "USGS:390735084333300:00011:00012",
  "USGS:390735084333300:00011:00013",
  "USGS:390735084333301:00011:00002",
  "USGS:390735084333301:00011:00001",
  "USGS:390735084333301:00011:00006",
  "USGS:09146200:00011:00001",
  "USGS:09146200:00011:00002",
  "USGS:09147000:00011:00015",
  "USGS:09147000:00011:00001",
  "USGS:09147000:00011:00002",
  "USGS:09147022:00011:00002",
  "USGS:09147022:00011:00001",
  "USGS:09147025:00011:00013",
  "USGS:09147025:00011:00011",
  "USGS:09147025:00011:00010",
  "USGS:09147500:00011:00017",
  "USGS:09147500:00011:00003",
  "USGS:09147500:00011:00001",
  "USGS:09147500:00011:00002",
  "USGS:09147500:00011:00019",
  "USGS:09149500:00011:00017",
  "USGS:09149500:00011:00001",
  "USGS:09149500:00011:00006",
  "USGS:09149500:00011:00019",
  "USGS:09152500:00011:00019",
  "USGS:09152500:00011:00001",
  "USGS:09152500:00011:00003",
  "USGS:09152500:00011:00020",
  "USGS:09163500:00011:00017",
  "USGS:09163500:00011:00001",
  "USGS:09163500:00011:00002",
  "USGS:09163500:00011:00018",
  "USGS:09165000:00011:00006",
  "USGS:09165000:00011:00004",
  "USGS:09166500:00011:00001",
  "USGS:09166500:00011:00002",
  "USGS:09166950:00011:00001",
  "USGS:09166950:00011:00002",
  "USGS:09168730:00011:00001",
  "USGS:09168730:00011:00002",
  "USGS:09169500:00011:00007",
  "USGS:09169500:00011:00006",
  "USGS:09169500:00011:00005",
  "USGS:09169500:00011:00008",
  "USGS:09171100:00011:00019",
  "USGS:09171100:00011:00001",
  "USGS:09171100:00011:00002",
  "USGS:09171100:00011:00020",
  "USGS:09171240:00011:00002",
  "USGS:09171240:00011:00001",
  "USGS:09171310:00011:00002",
  "USGS:09171310:00011:00001",
  "USGS:09172500:00011:00001",
  "USGS:09172500:00011:00004",
  "USGS:09174600:00011:00002",
  "USGS:09174600:00011:00001",
  "USGS:09177000:00011:00001",
  "USGS:09177000:00011:00002",
  "USGS:09179450:00011:00001",
  "USGS:09237450:00011:00002",
  "USGS:09237450:00011:00003",
  "USGS:09237500:00011:00002",
  "USGS:09237500:00011:00001",
  "USGS:09238900:00011:00001",
  "USGS:09238900:00011:00003",
  "USGS:09239500:00011:00004",
  "USGS:09239500:00011:00003",
  "USGS:09240020:00011:00001",
  "USGS:09240020:00011:00002",
  "USGS:09242500:00011:00001",
  "USGS:09242500:00011:00004",
  "USGS:09244490:00011:00002",
  "USGS:09244490:00011:00001",
  "USGS:09246200:00011:00001",
  "USGS:09246200:00011:00002",
  "USGS:09246500:00011:00001",
  "USGS:09246500:00011:00002",
  "USGS:09247600:00011:00001",
  "USGS:09247600:00011:00003",
  "USGS:09251000:00011:00005",
  "USGS:09251000:00011:00001",
  "USGS:09251000:00011:00002",
  "USGS:09251000:00011:00016",
  "USGS:09251000:00011:00026",
  "USGS:09253000:00011:00004",
  "USGS:09253000:00011:00002",
  "USGS:09255000:00011:00001",
  "USGS:09255000:00011:00004",
  "USGS:09260000:00011:00006",
  "USGS:09260000:00011:00002",
  "USGS:09260050:00011:00001",
  "USGS:09260050:00011:00006",
  "USGS:09260050:00011:00005",
  "USGS:09304200:00011:00001",
  "USGS:09304200:00011:00002",
  "USGS:09304200:00011:00006",
  "USGS:09304500:00011:00003",
  "USGS:09304500:00011:00005",
  "USGS:09304800:00011:00001",
  "USGS:09304800:00011:00002",
  "USGS:09304800:00011:00006",
  "USGS:09304800:00011:00003",
  "USGS:09306200:00011:00008",
  "USGS:09306200:00011:00002",
  "USGS:09306200:00011:00007",
  "USGS:09306200:00011:00009",
  "USGS:09306222:00011:00001",
  "USGS:09306222:00011:00003",
  "USGS:09306222:00011:00008",
  "USGS:09306222:00011:00004",
  "USGS:09306242:00011:00002",
  "USGS:09306242:00011:00007",
  "USGS:09306255:00011:00001",
  "USGS:09306255:00011:00003",
  "USGS:09306255:00011:00008",
  "USGS:09306255:00011:00004",
  "USGS:09306290:00011:00015",
  "USGS:09306290:00011:00001",
  "USGS:09306290:00011:00002",
  "USGS:09306290:00011:00016",
  "USGS:09342500:00011:00001",
  "USGS:09342500:00011:00002",
  "USGS:09346400:00011:00001",
  "USGS:09346400:00011:00003",
  "USGS:09349800:00011:00001",
  "USGS:09349800:00011:00002",
  "USGS:09352900:00011:00002",
  "USGS:09352900:00011:00001",
  "USGS:01377000:00011:00001",
  "USGS:01377000:00011:00002",
  "USGS:01377370:00011:00002",
  "USGS:01377370:00011:00001",
  "USGS:01377450:00011:00001",
  "USGS:01377451:00011:00013",
  "USGS:01377451:00011:00001",
  "USGS:01377500:00011:00001",
  "USGS:01377500:00011:00002",
  "USGS:01378480:00011:00001",
  "USGS:01378500:00011:00001",
  "USGS:01378500:00011:00002",
  "USGS:01379000:00011:00001",
  "USGS:01379000:00011:00002",
  "USGS:01379500:00011:00002",
  "USGS:01379500:00011:00005",
  "USGS:01379530:00011:00009",
  "USGS:01379530:00011:00001",
  "USGS:01379530:00011:00002",
  "USGS:01379530:00011:00004",
  "USGS:01379699:00011:00002",
  "USGS:01379699:00011:00001",
  "USGS:01379773:00011:00002",
  "USGS:01379773:00011:00006",
  "USGS:01379780:00011:00001",
  "USGS:01379780:00011:00002",
  "USGS:01379845:00011:00001",
  "USGS:07152000:00011:00015",
  "USGS:07152000:00011:00007",
  "USGS:07152000:00011:00006",
  "USGS:07152500:00011:00013",
  "USGS:07152500:00011:00012",
  "USGS:07153000:00011:00014",
  "USGS:07153000:00011:00004",
  "USGS:07153000:00011:00015",
  "USGS:07154500:00011:00006",
  "USGS:07154500:00011:00005",
  "USGS:07154500:00011:00004",
  "USGS:07157950:00011:00014",
  "USGS:07157950:00011:00013",
  "USGS:07157950:00011:00012",
  "USGS:07158000:00011:00023",
  "USGS:07158000:00011:00013",
  "USGS:07158000:00011:00012",
  "USGS:07159100:00011:00012",
  "USGS:07159100:00011:00011",
  "USGS:07159550:00011:00015",
  "USGS:07159550:00011:00002",
  "USGS:07159550:00011:00001",
  "USGS:07159550:00011:00014",
  "USGS:07159750:00011:00016",
  "USGS:07159750:00011:00018",
  "USGS:07159750:00011:00017",
  "USGS:07160000:00011:00005",
  "USGS:07160000:00011:00004",
  "USGS:07160000:00011:00015",
  "USGS:07160350:00011:00014",
  "USGS:07160350:00011:00003",
  "USGS:07160350:00011:00002",
  "USGS:07160350:00011:00001",
  "USGS:07160350:00011:00015",
  "USGS:385117107554501:00011:00001",
  "USGS:385121104480701:00011:00002",
  "USGS:385129104544601:00011:00002",
  "USGS:385240104444801:00011:00002",
  "USGS:385241104560101:00011:00002",
  "USGS:385259104410801:00011:00002",
  "USGS:385334104544901:00011:00002",
  "USGS:385349104501401:00011:00002",
  "USGS:385449104565501:00011:00002",
  "USGS:385519104415501:00011:00002",
  "USGS:385520104530401:00011:00002",
  "USGS:385548104503201:00011:00002",
  "USGS:385636104465601:00011:00002",
  "USGS:385740104405501:00011:00002",
  "USGS:385846104462501:00011:00002",
  "USGS:385906104495101:00011:00002",
  "USGS:391517106223801:00011:00002",
  "USGS:391517106223801:00011:00001",
  "USGS:393109104464500:00011:00002",
  "USGS:393109104464500:00011:00003",
  "USGS:393803107435601:00011:00001",
  "USGS:393839107463801:00011:00001",
  "USGS:393938104572101:00011:00002",
  "USGS:393947104555101:00011:00002",
  "USGS:394028104560201:00011:00002",
  "USGS:394028104565501:00011:00002",
  "USGS:394220106431500:00011:00003",
  "USGS:394220106431500:00011:00002",
  "USGS:394220106431500:00011:00001",
  "USGS:394220106431500:00011:00004",
  "USGS:394308105413800:00011:00002",
  "USGS:394308105413800:00011:00001",
  "USGS:394329104490101:00011:00002",
  "USGS:394329104490101:00011:00001",
  "USGS:394359105411901:00011:00001",
  "USGS:394839104570300:00011:00002",
  "USGS:394839104570300:00011:00021",
  "USGS:401638105402601:00011:00003",
  "USGS:401719105394311:00011:00003",
  "USGS:401719105394311:00011:00006",
  "USGS:401723105400101:00011:00006",
  "USGS:401733105392404:00011:00007",
  "USGS:402114105350101:00011:00015",
  "USGS:402114105350101:00011:00002",
  "USGS:402114105350101:00011:00003",
  "USGS:402214104255101:00011:00002",
  "USGS:402214104255101:00011:00001",
  "USGS:404417108524900:00011:00001",
  "USGS:01383500:00011:00001",
  "USGS:01383500:00011:00002",
  "USGS:03136500:00011:00004",
  "USGS:03136500:00011:00003",
  "USGS:03138500:00011:00004",
  "USGS:03139000:00011:00007",
  "USGS:03139000:00011:00006",
  "USGS:03139850:00011:00001",
  "USGS:03140000:00011:00001",
  "USGS:03140000:00011:00002",
  "USGS:03140500:00011:00004",
  "USGS:03140500:00011:00003",
  "USGS:03141500:00011:00003",
  "USGS:03141700:00011:00001",
  "USGS:03141870:00011:00002",
  "USGS:03141870:00011:00001",
  "USGS:03142000:00011:00006",
  "USGS:03142000:00011:00005",
  "USGS:03143500:00011:00003",
  "USGS:03144000:00011:00004",
  "USGS:03144000:00011:00003",
  "USGS:03144500:00011:00002",
  "USGS:03144500:00011:00006",
  "USGS:03144816:00011:00003",
  "USGS:03144816:00011:00002",
  "USGS:03144816:00011:00001",
  "USGS:03144950:00011:00001",
  "USGS:03145000:00011:00004",
  "USGS:03145000:00011:00003",
  "USGS:03145173:00011:00011",
  "USGS:03145173:00011:00001",
  "USGS:03145483:00011:00003",
  "USGS:03145483:00011:00002",
  "USGS:03145483:00011:00001",
  "USGS:03145534:00011:00002",
  "USGS:03145534:00011:00001",
  "USGS:03146000:00011:00002",
  "USGS:03146000:00011:00003",
  "USGS:03146277:00011:00012",
  "USGS:03146277:00011:00001",
  "USGS:03146402:00011:00011",
  "USGS:03146402:00011:00001",
  "USGS:03146405:00011:00003",
  "USGS:03146405:00011:00001",
  "USGS:03146500:00011:00010",
  "USGS:03146500:00011:00009",
  "USGS:03147500:00011:00001",
  "USGS:03148000:00011:00003",
  "USGS:03149500:00011:00001",
  "USGS:03149500:00011:00002",
  "USGS:03150000:00011:00002",
  "USGS:03150000:00011:00001",
  "USGS:03150500:00011:00011",
  "USGS:03150500:00011:00001",
  "USGS:03150700:00011:00002",
  "USGS:03150700:00011:00001",
  "USGS:03157000:00011:00004",
  "USGS:03157000:00011:00001",
  "USGS:03157000:00011:00002",
  "USGS:03157500:00011:00004",
  "USGS:03157500:00011:00003",
  "USGS:03158200:00011:00004",
  "USGS:03158510:00011:00001",
  "USGS:03159000:00011:00003",
  "USGS:03159246:00011:00002",
  "USGS:03159246:00011:00001",
  "USGS:03159500:00011:00008",
  "USGS:03159500:00011:00007",
  "USGS:03159540:00011:00016",
  "USGS:03159540:00011:00004",
  "USGS:03159540:00011:00003",
  "USGS:03201902:00011:00001",
  "USGS:03201902:00011:00004",
  "USGS:03201980:00011:00006",
  "USGS:03201980:00011:00005",
  "USGS:03202000:00011:00010",
  "USGS:03202000:00011:00009",
  "USGS:01398500:00011:00002",
  "USGS:01398500:00011:00003",
  "USGS:01398900:00011:00002",
  "USGS:01398900:00011:00001",
  "USGS:01399100:00011:00001",
  "USGS:01399100:00011:00002",
  "USGS:01399100:00011:00003",
  "USGS:01399500:00011:00001",
  "USGS:01399500:00011:00002",
  "USGS:01399670:00011:00001",
  "USGS:01399670:00011:00002",
  "USGS:01399780:00011:00001",
  "USGS:01399830:00011:00002",
  "USGS:01400000:00011:00001",
  "USGS:01400000:00011:00002",
  "USGS:03221500:00011:00003",
  "USGS:03221500:00011:00004",
  "USGS:03221500:00011:00005",
  "USGS:03221500:00011:00006",
  "USGS:03221500:00011:00002",
  "USGS:03221646:00011:00001",
  "USGS:03223000:00011:00003",
  "USGS:03223425:00011:00002",
  "USGS:03223425:00011:00001",
  "USGS:03225500:00011:00005",
  "USGS:03225500:00011:00004",
  "USGS:03226800:00011:00016",
  "USGS:03226800:00011:00001",
  "USGS:03227500:00011:00001",
  "USGS:03227500:00011:00002",
  "USGS:03228039:00011:00001",
  "USGS:03228039:00011:00002",
  "USGS:03228039:00011:00003",
  "USGS:03228039:00011:00004",
  "USGS:03228039:00011:00005",
  "USGS:03228300:00011:00005",
  "USGS:03228300:00011:00004",
  "USGS:03228300:00011:00003",
  "USGS:03228300:00011:00006",
  "USGS:03228300:00011:00007",
  "USGS:03228300:00011:00008",
  "USGS:03228400:00011:00002",
  "USGS:03228500:00011:00004",
  "USGS:03228500:00011:00003",
  "USGS:03228750:00011:00012",
  "USGS:03228750:00011:00001",
  "USGS:03228805:00011:00008",
  "USGS:03228805:00011:00006",
  "USGS:03228805:00011:00005",
  "USGS:03229000:00011:00001",
  "USGS:03229500:00011:00004",
  "USGS:03229500:00011:00003",
  "USGS:03229610:00011:00002",
  "USGS:03229610:00011:00001",
  "USGS:03229796:00011:00002",
  "USGS:03229796:00011:00001",
  "USGS:03230310:00011:00017",
  "USGS:03230310:00011:00002",
  "USGS:03230310:00011:00001",
  "USGS:03230450:00011:00002",
  "USGS:03230450:00011:00001",
  "USGS:03230500:00011:00004",
  "USGS:03230500:00011:00003",
  "USGS:03230700:00011:00001",
  "USGS:03230700:00011:00003",
  "USGS:03230800:00011:00015",
  "USGS:03230800:00011:00003",
  "USGS:03230900:00011:00003",
  "USGS:03231000:00011:00005",
  "USGS:03231500:00011:00036",
  "USGS:03231500:00011:00008",
  "USGS:03231500:00011:00007",
  "USGS:03232000:00011:00016",
  "USGS:03232000:00011:00005",
  "USGS:03232300:00011:00003",
  "USGS:03232470:00011:00006",
  "USGS:03232470:00011:00003",
  "USGS:03232500:00011:00004",
  "USGS:03232500:00011:00003",
  "USGS:03234000:00011:00021",
  "USGS:03234000:00011:00002",
  "USGS:03234000:00011:00007",
  "USGS:03234300:00011:00014",
  "USGS:03234300:00011:00013",
  "USGS:03234500:00011:00002",
  "USGS:03234500:00011:00001",
  "USGS:03237020:00011:00002",
  "USGS:03237020:00011:00003",
  "USGS:03237280:00011:00016",
  "USGS:03237280:00011:00015",
  "USGS:03237500:00011:00015",
  "USGS:03237500:00011:00001",
  "USGS:03237500:00011:00002",
  "USGS:03238495:00011:00002",
  "USGS:03238495:00011:00001",
  "USGS:03240000:00011:00001",
  "USGS:03240000:00011:00002",
  "USGS:03240000:00011:00005",
  "USGS:03241500:00011:00003",
  "USGS:03241500:00011:00001",
  "USGS:03242050:00011:00007",
  "USGS:03242340:00011:00001",
  "USGS:03242340:00011:00002",
  "USGS:03242350:00011:00005",
  "USGS:03242350:00011:00003",
  "USGS:03244936:00011:00002",
  "USGS:03244936:00011:00001",
  "USGS:01409334:00011:00004",
  "USGS:01409334:00011:00002",
  "USGS:01409334:00011:00001",
  "USGS:01409335:00011:00005",
  "USGS:01409335:00011:00001",
  "USGS:01409400:00011:00001",
  "USGS:01409400:00011:00013",
  "USGS:01409810:00011:00002",
  "USGS:01409810:00011:00014",
  "USGS:01410000:00011:00001",
  "USGS:01410000:00011:00002",
  "USGS:01410150:00011:00001",
  "USGS:01410150:00011:00002",
  "USGS:01410500:00011:00002",
  "USGS:01410500:00011:00003",
  "USGS:01410510:00011:00005",
  "USGS:01410510:00011:00001",
  "USGS:01410560:00011:00015",
  "USGS:01410560:00011:00001",
  "USGS:01410600:00011:00016",
  "USGS:01410600:00011:00001",
  "USGS:01410784:00011:00002",
  "USGS:01410784:00011:00001",
  "USGS:01410820:00011:00001",
  "USGS:01410820:00011:00002",
  "USGS:01411000:00011:00003",
  "USGS:01411000:00011:00007",
  "USGS:01411300:00011:00014",
  "USGS:01411300:00011:00001",
  "USGS:390735084333301:00011:00007",
  "USGS:390735084333301:00011:00008",
  "USGS:390841082535800:00011:00001",
  "USGS:390844084322201:00011:00001",
  "USGS:390844084322202:00011:00001",
  "USGS:391214084470100:00011:00003",
  "USGS:391214084470100:00011:00002",
  "USGS:391905084381000:00011:00001",
  "USGS:392016082272400:00011:00001",
  "USGS:392236084334800:00011:00001",
  "USGS:392553081281600:00011:00002",
  "USGS:392808084283600:00011:00001",
  "USGS:392902084255900:00011:00001",
  "USGS:393153083322000:00011:00001",
  "USGS:393318084190100:00011:00001",
  "USGS:394442084111600:00011:00001",
  "USGS:394533084113800:00011:00002",
  "USGS:394533084113800:00011:00001",
  "USGS:394915084103300:00011:00001",
  "USGS:395316083593100:00011:00001",
  "USGS:395417082314200:00011:00003",
  "USGS:395417082314200:00011:00015",
  "USGS:395417082314200:00011:00004",
  "USGS:395417082314200:00011:00014",
  "USGS:395521081260500:00011:00007",
  "USGS:395521081260500:00011:00003",
  "USGS:395521081260500:00011:00004",
  "USGS:395521081260500:00011:00001",
  "USGS:395521081260500:00011:00005",
  "USGS:395521081260500:00011:00009",
  "USGS:395521081260500:00011:00006",
  "USGS:395521081260500:00011:00008",
  "USGS:395847084085500:00011:00002",
  "USGS:395847084085500:00011:00001",
  "USGS:400150083053401:00011:00002",
  "USGS:400150083053401:00011:00001",
  "USGS:400150083053402:00011:00002",
  "USGS:400150083053402:00011:00001",
  "USGS:400151083053400:00011:00007",
  "USGS:400151083053400:00011:00003",
  "USGS:400151083053400:00011:00004",
  "USGS:400151083053400:00011:00001",
  "USGS:400151083053400:00011:00005",
  "USGS:400151083053400:00011:00008",
  "USGS:400151083053400:00011:00009",
  "USGS:400153083053600:00011:00002",
  "USGS:400153083053600:00011:00001",
  "USGS:400540082540400:00011:00003",
  "USGS:401122084143400:00011:00001",
  "USGS:401133081125300:00011:00007",
  "USGS:401133081125300:00011:00003",
  "USGS:401133081125300:00011:00004",
  "USGS:401133081125300:00011:00001",
  "USGS:401133081125300:00011:00005",
  "USGS:401133081125300:00011:00009",
  "USGS:401133081125300:00011:00006",
  "USGS:03255420:00011:00001",
  "USGS:401133081125300:00011:00008",
  "USGS:402120081134200:00011:00007",
  "USGS:402120081134200:00011:00003",
  "USGS:402120081134200:00011:00004",
  "USGS:402120081134200:00011:00001",
  "USGS:402120081134200:00011:00005",
  "USGS:402120081134200:00011:00009",
  "USGS:402120081134200:00011:00006",
  "USGS:402120081134200:00011:00008",
  "USGS:402815081114300:00011:00007",
  "USGS:402815081114300:00011:00003",
  "USGS:402815081114300:00011:00004",
  "USGS:402815081114300:00011:00001",
  "USGS:402815081114300:00011:00005",
  "USGS:402815081114300:00011:00009",
  "USGS:402815081114300:00011:00006",
  "USGS:402815081114300:00011:00008",
  "USGS:402913084285400:00011:00002",
  "USGS:402913084285400:00011:00001",
  "USGS:402913084285400:00011:00003",
  "USGS:402958084363300:00011:00018",
  "USGS:402958084363300:00011:00002",
  "USGS:402958084363300:00011:00001",
  "USGS:403127081171000:00011:00007",
  "USGS:403127081171000:00011:00003",
  "USGS:403127081171000:00011:00004",
  "USGS:403127081171000:00011:00001",
  "USGS:403127081171000:00011:00005",
  "USGS:403127081171000:00011:00009",
  "USGS:403127081171000:00011:00006",
  "USGS:403127081171000:00011:00008",
  "USGS:404648083412600:00011:00002",
  "USGS:404655081553100:00011:00002",
  "USGS:405051083391001:00011:00002",
  "USGS:405051083391001:00011:00001",
  "USGS:405051083391001:00011:00005",
  "USGS:410014081362600:00011:00018",
  "USGS:410014081362600:00011:00002",
  "USGS:410014081362600:00011:00001",
  "USGS:410121081330300:00011:00003",
  "USGS:410121081330300:00011:00001",
  "USGS:410433081312500:00011:00002",
  "USGS:410433081312500:00011:00001",
  "USGS:411438081085200:00011:00001",
  "USGS:411819082493900:00011:00001",
  "USGS:412141081412100:00011:00002",
  "USGS:412141081412100:00011:00001",
  "USGS:412325081415500:00011:00002",
  "USGS:412325081415500:00011:00001",
  "USGS:412453081395500:00011:00011",
  "USGS:412453081395500:00011:00001",
  "USGS:412533081221500:00011:00002",
  "USGS:412533081221500:00011:00001",
  "USGS:412624081450700:00011:00002",
  "USGS:412624081450700:00011:00001",
  "USGS:01463620:00011:00001",
  "USGS:03255500:00011:00002",
  "USGS:03256500:00011:00001",
  "USGS:03259000:00011:00001",
  "USGS:03259000:00011:00002",
  "USGS:03259973:00011:00002",
  "USGS:03259973:00011:00001",
  "USGS:03260706:00011:00006",
  "USGS:03260706:00011:00005",
  "USGS:03260706:00011:00004",
  "USGS:03260706:00011:00007",
  "USGS:03261500:00011:00019",
  "USGS:03261500:00011:00008",
  "USGS:03261500:00011:00002",
  "USGS:03261500:00011:00005",
  "USGS:03261500:00011:00010",
  "USGS:03261950:00011:00002",
  "USGS:03261950:00011:00003",
  "USGS:03261950:00011:00006",
  "USGS:03261950:00011:00010",
  "USGS:03262000:00011:00001",
  "USGS:03262000:00011:00002",
  "USGS:03262000:00011:00004",
  "USGS:03262500:00011:00001",
  "USGS:03262500:00011:00002",
  "USGS:03262500:00011:00003",
  "USGS:03262700:00011:00001",
  "USGS:03262700:00011:00002",
  "USGS:03262700:00011:00004",
  "USGS:03263000:00011:00005",
  "USGS:03263000:00011:00001",
  "USGS:03263000:00011:00002",
  "USGS:03263000:00011:00007",
  "USGS:03264000:00011:00001",
  "USGS:03264000:00011:00002",
  "USGS:03264000:00011:00004",
  "USGS:03265000:00011:00004",
  "USGS:03265000:00011:00003",
  "USGS:03265000:00011:00001",
  "USGS:03265000:00011:00006",
  "USGS:03266000:00011:00004",
  "USGS:03266000:00011:00001",
  "USGS:03266000:00011:00002",
  "USGS:03266000:00011:00005",
  "USGS:03266560:00011:00002",
  "USGS:03266560:00011:00001",
  "USGS:03267000:00011:00005",
  "USGS:03267000:00011:00004",
  "USGS:03267000:00011:00003",
  "USGS:03267000:00011:00008",
  "USGS:03267900:00011:00014",
  "USGS:03267900:00011:00004",
  "USGS:03267900:00011:00003",
  "USGS:03267900:00011:00005",
  "USGS:03268090:00011:00001",
  "USGS:03269500:00011:00014",
  "USGS:03269500:00011:00001",
  "USGS:03269500:00011:00002",
  "USGS:03269500:00011:00015",
  "USGS:03270000:00011:00012",
  "USGS:03270000:00011:00003",
  "USGS:03270000:00011:00008",
  "USGS:03270000:00011:00014",
  "USGS:03270500:00011:00003",
  "USGS:03270500:00011:00002",
  "USGS:03270500:00011:00005",
  "USGS:03271000:00011:00001",
  "USGS:03271000:00011:00002",
  "USGS:03271000:00011:00004",
  "USGS:03271207:00011:00001",
  "USGS:03271207:00011:00002",
  "USGS:03271300:00011:00002",
  "USGS:03271300:00011:00001",
  "USGS:03271300:00011:00007",
  "USGS:03271500:00011:00001",
  "USGS:03271500:00011:00006",
  "USGS:03271601:00011:00014",
  "USGS:03271601:00011:00002",
  "USGS:03271601:00011:00001",
  "USGS:03271620:00011:00011",
  "USGS:03271620:00011:00001",
  "USGS:03271620:00011:00002",
  "USGS:03272000:00011:00013",
  "USGS:03272000:00011:00001",
  "USGS:03272000:00011:00002",
  "USGS:03272000:00011:00004",
  "USGS:03272100:00011:00003",
  "USGS:03272100:00011:00002",
  "USGS:03272100:00011:00001",
  "USGS:03272100:00011:00004",
  "USGS:03272700:00011:00005",
  "USGS:03272700:00011:00001",
  "USGS:03272700:00011:00002",
  "USGS:03272700:00011:00007",
  "USGS:03274000:00011:00003",
  "USGS:03274000:00011:00001",
  "USGS:03274000:00011:00002",
  "USGS:03274000:00011:00007",
  "USGS:03274615:00011:00001",
  "USGS:03322485:00011:00001",
  "USGS:04177000:00011:00004",
  "USGS:04177000:00011:00003",
  "USGS:04178000:00011:00001",
  "USGS:04178000:00011:00004",
  "USGS:04180988:00011:00004",
  "USGS:04180988:00011:00003",
  "USGS:04180988:00011:00002",
  "USGS:04180988:00011:00001",
  "USGS:04183500:00011:00003",
  "USGS:04183500:00011:00004",
  "USGS:04183500:00011:00005",
  "USGS:04184500:00011:00001",
  "USGS:04184500:00011:00004",
  "USGS:04185000:00011:00015",
  "USGS:04185000:00011:00004",
  "USGS:04185000:00011:00003",
  "USGS:04185318:00011:00001",
  "USGS:04185318:00011:00002",
  "USGS:394652075100401:00011:00001",
  "USGS:394652075100402:00011:00001",
  "USGS:394728074452501:00011:00001",
  "USGS:394800074524601:00011:00001",
  "USGS:03090500:00011:00003",
  "USGS:03091000:00011:00011",
  "USGS:03091000:00011:00015",
  "USGS:03091500:00011:00014",
  "USGS:03091500:00011:00004",
  "USGS:03091500:00011:00003",
  "USGS:03092090:00011:00015",
  "USGS:03092090:00011:00003",
  "USGS:03092090:00011:00001",
  "USGS:03092450:00011:00013",
  "USGS:03092460:00011:00015",
  "USGS:03092460:00011:00005",
  "USGS:03092460:00011:00004",
  "USGS:03092460:00011:00003",
  "USGS:03093000:00011:00004",
  "USGS:03093000:00011:00003",
  "USGS:03094000:00011:00015",
  "USGS:03094000:00011:00014",
  "USGS:03094000:00011:00003",
  "USGS:03094000:00011:00001",
  "USGS:03094704:00011:00002",
  "USGS:03094704:00011:00012",
  "USGS:03094704:00011:00001",
  "USGS:03095000:00011:00012",
  "USGS:03095500:00011:00015",
  "USGS:03095500:00011:00005",
  "USGS:03095500:00011:00004",
  "USGS:03095500:00011:00001",
  "USGS:03098600:00011:00016",
  "USGS:03098600:00011:00025",
  "USGS:03098600:00011:00002",
  "USGS:03098600:00011:00001",
  "USGS:03098600:00011:00018",
  "USGS:03098600:00011:00019",
  "USGS:03098600:00011:00017",
  "USGS:03098700:00011:00002",
  "USGS:03098700:00011:00001",
  "USGS:03099500:00011:00019",
  "USGS:03099500:00011:00008",
  "USGS:03099500:00011:00007",
  "USGS:03099500:00011:00003",
  "USGS:03102950:00011:00016",
  "USGS:03102950:00011:00014",
  "USGS:03102950:00011:00001",
  "USGS:03109500:00011:00001",
  "USGS:03109500:00011:00002",
  "USGS:03110000:00011:00004",
  "USGS:03110000:00011:00003",
  "USGS:03110685:00011:00001",
  "USGS:03110690:00011:00002",
  "USGS:03110690:00011:00001",
  "USGS:03111500:00011:00004",
  "USGS:03111500:00011:00001",
  "USGS:03111548:00011:00019",
  "USGS:03111548:00011:00006",
  "USGS:03111548:00011:00005",
  "USGS:03113990:00011:00002",
  "USGS:03113990:00011:00001",
  "USGS:03114275:00011:00001",
  "USGS:03114280:00011:00012",
  "USGS:03114280:00011:00001",
  "USGS:03114306:00011:00002",
  "USGS:03114306:00011:00003",
  "USGS:03114306:00011:00001",
  "USGS:03115400:00011:00004",
  "USGS:03115400:00011:00003",
  "USGS:03115644:00011:00002",
  "USGS:03115644:00011:00001",
  "USGS:03115712:00011:00003",
  "USGS:03115712:00011:00002",
  "USGS:03115712:00011:00001",
  "USGS:03115786:00011:00002",
  "USGS:03115786:00011:00001",
  "USGS:03115973:00011:00002",
  "USGS:03115973:00011:00001",
  "USGS:03116077:00011:00013",
  "USGS:03116077:00011:00002",
  "USGS:03116077:00011:00003",
  "USGS:03117000:00011:00004",
  "USGS:03117000:00011:00003",
  "USGS:03117500:00011:00004",
  "USGS:03117500:00011:00003",
  "USGS:03118000:00011:00004",
  "USGS:03118000:00011:00003",
  "USGS:03118500:00011:00004",
  "USGS:03118500:00011:00003",
  "USGS:03120500:00011:00005",
  "USGS:03120500:00011:00003",
  "USGS:03121500:00011:00002",
  "USGS:03121850:00011:00006",
  "USGS:03121850:00011:00004",
  "USGS:03121850:00011:00003",
  "USGS:03121850:00011:00008",
  "USGS:03121850:00011:00010",
  "USGS:03121850:00011:00012",
  "USGS:03122500:00011:00003",
  "USGS:03124000:00011:00003",
  "USGS:03124500:00011:00001",
  "USGS:03124500:00011:00002",
  "USGS:03124800:00011:00012",
  "USGS:03124800:00011:00001",
  "USGS:03125900:00011:00001",
  "USGS:03126000:00011:00003",
  "USGS:03126910:00011:00003",
  "USGS:03126910:00011:00001",
  "USGS:07160500:00011:00006",
  "USGS:07160500:00011:00005",
  "USGS:07160500:00011:00004",
  "USGS:07160810:00011:00001",
  "USGS:402805074385601:00011:00001",
  "USGS:402955074312501:00011:00001",
  "USGS:403200074420601:00011:00001",
  "USGS:403300074202901:00011:00001",
  "USGS:403328074434901:00011:00001",
  "USGS:403338074325301:00011:00001",
  "USGS:403430074365701:00011:00001",
  "USGS:403455074514801:00011:00001",
  "USGS:403506074302801:00011:00001",
  "USGS:403517074452501:00011:00001",
  "USGS:01400010:00011:00001",
  "USGS:01400360:00011:00001",
  "USGS:01400500:00011:00018",
  "USGS:01400500:00011:00001",
  "USGS:01400500:00011:00002",
  "USGS:01400500:00011:00020",
  "USGS:01400500:00011:00022",
  "USGS:01400500:00011:00021",
  "USGS:01400500:00011:00019",
  "USGS:01400500:00011:00023",
  "USGS:01401000:00011:00002",
  "USGS:01401000:00011:00005",
  "USGS:01401650:00011:00002",
  "USGS:01401650:00011:00003",
  "USGS:01401750:00011:00013",
  "USGS:01401750:00011:00001",
  "USGS:01402000:00011:00001",
  "USGS:01402000:00011:00002",
  "USGS:01402500:00011:00004",
  "USGS:01402500:00011:00001",
  "USGS:01402540:00011:00012",
  "USGS:01402540:00011:00001",
  "USGS:01402630:00011:00001",
  "USGS:01402630:00011:00002",
  "USGS:01403060:00011:00001",
  "USGS:01403060:00011:00002",
  "USGS:01403150:00011:00002",
  "USGS:01403150:00011:00003",
  "USGS:01403200:00011:00001",
  "USGS:01403400:00011:00002",
  "USGS:01403400:00011:00003",
  "USGS:01403540:00011:00001",
  "USGS:01403540:00011:00002",
  "USGS:01403570:00011:00001",
  "USGS:01403600:00011:00001",
  "USGS:01403900:00011:00005",
  "USGS:01403900:00011:00004",
  "USGS:01405030:00011:00002",
  "USGS:01405030:00011:00001",
  "USGS:01405400:00011:00001",
  "USGS:01405400:00011:00002",
  "USGS:01406050:00011:00002",
  "USGS:01406050:00011:00001",
  "USGS:01406710:00011:00004",
  "USGS:01406710:00011:00001",
  "USGS:01407081:00011:00019",
  "USGS:01407081:00011:00001",
  "USGS:01407290:00011:00002",
  "USGS:01407290:00011:00012",
  "USGS:01407498:00011:00001",
  "USGS:01407498:00011:00002",
  "USGS:01407500:00011:00001",
  "USGS:01407500:00011:00002",
  "USGS:01407600:00011:00005",
  "USGS:01407600:00011:00001",
  "USGS:01407705:00011:00001",
  "USGS:01407705:00011:00002",
  "USGS:01407760:00011:00001",
  "USGS:01407760:00011:00002",
  "USGS:01407770:00011:00003",
  "USGS:01407770:00011:00001",
  "USGS:01408000:00011:00001",
  "USGS:01408000:00011:00002",
  "USGS:01408000:00011:00006",
  "USGS:01408000:00011:00003",
  "USGS:01408000:00011:00018",
  "USGS:01408029:00011:00013",
  "USGS:01408029:00011:00002",
  "USGS:01408029:00011:00001",
  "USGS:01408029:00011:00014",
  "USGS:01408029:00011:00015",
  "USGS:01408048:00011:00003",
  "USGS:01408048:00011:00001",
  "USGS:01408120:00011:00001",
  "USGS:01408120:00011:00002",
  "USGS:01408168:00011:00007",
  "USGS:01408168:00011:00002",
  "USGS:01408205:00011:00004",
  "USGS:01408205:00011:00002",
  "USGS:01408205:00011:00001",
  "USGS:01408500:00011:00001",
  "USGS:01408500:00011:00002",
  "USGS:01408500:00011:00005",
  "USGS:01408500:00011:00003",
  "USGS:01408500:00011:00018",
  "USGS:01408500:00011:00017",
  "USGS:01408500:00011:00004",
  "USGS:01408500:00011:00016",
  "USGS:01408500:00011:00021",
  "USGS:01408900:00011:00002",
  "USGS:01408900:00011:00001",
  "USGS:01409125:00011:00019",
  "USGS:01409125:00011:00001",
  "USGS:01409146:00011:00015",
  "USGS:01409146:00011:00020",
  "USGS:01409146:00011:00019",
  "USGS:01409147:00011:00004",
  "USGS:01409147:00011:00002",
  "USGS:01409147:00011:00001",
  "USGS:01409280:00011:00013",
  "USGS:01409280:00011:00001",
  "USGS:01409280:00011:00002",
  "USGS:01427207:00011:00015",
  "USGS:01427207:00011:00012",
  "USGS:01427207:00011:00004",
  "USGS:01427510:00011:00003",
  "USGS:01427510:00011:00007",
  "USGS:01427510:00011:00002",
  "USGS:01427510:00011:00005",
  "USGS:01428750:00011:00006",
  "USGS:01428750:00011:00005",
  "USGS:01428750:00011:00004",
  "USGS:01428750:00011:00003",
  "USGS:01428900:00011:00001",
  "USGS:01429000:00011:00003",
  "USGS:01429000:00011:00013",
  "USGS:01429000:00011:00001",
  "USGS:01429000:00011:00002",
  "USGS:01429400:00011:00001",
  "USGS:01429500:00011:00012",
  "USGS:01379868:00011:00003",
  "USGS:01379868:00011:00002",
  "USGS:01379868:00011:00001",
  "USGS:01380450:00011:00002",
  "USGS:01380450:00011:00001",
  "USGS:01380900:00011:00002",
  "USGS:01381000:00011:00001",
  "USGS:01381000:00011:00002",
  "USGS:01381400:00011:00002",
  "USGS:01381400:00011:00001",
  "USGS:01381500:00011:00001",
  "USGS:01381500:00011:00002",
  "USGS:01381800:00011:00002",
  "USGS:01381800:00011:00001",
  "USGS:01381900:00011:00001",
  "USGS:01381900:00011:00002",
  "USGS:01381940:00011:00001",
  "USGS:01382170:00011:00012",
  "USGS:01382170:00011:00001",
  "USGS:01382170:00011:00002",
  "USGS:01382210:00011:00003",
  "USGS:01382210:00011:00002",
  "USGS:01382210:00011:00001",
  "USGS:01382210:00011:00005",
  "USGS:01382210:00011:00007",
  "USGS:01382210:00011:00006",
  "USGS:01382270:00011:00002",
  "USGS:01382270:00011:00001",
  "USGS:01382310:00011:00001",
  "USGS:01382381:00011:00001",
  "USGS:01382385:00011:00003",
  "USGS:01382385:00011:00002",
  "USGS:01382385:00011:00001",
  "USGS:01382500:00011:00014",
  "USGS:01382500:00011:00001",
  "USGS:01382500:00011:00002",
  "USGS:01382800:00011:00002",
  "USGS:01382800:00011:00001",
  "USGS:01383000:00011:00002",
  "USGS:10396000:00011:00013",
  "USGS:10396000:00011:00002",
  "USGS:10396000:00011:00001",
  "USGS:11486990:00011:00005",
  "USGS:11486990:00011:00010",
  "USGS:11486990:00011:00003",
  "USGS:11492200:00011:00003",
  "USGS:11493500:00011:00001",
  "USGS:11493500:00011:00002",
  "USGS:11497550:00011:00001",
  "USGS:11501000:00011:00003",
  "USGS:11501000:00011:00001",
  "USGS:11501000:00011:00002",
  "USGS:11501000:00011:00008",
  "USGS:11502500:00011:00010",
  "USGS:11502500:00011:00001",
  "USGS:11502500:00011:00002",
  "USGS:11502500:00011:00007",
  "USGS:11503000:00011:00001",
  "USGS:11503000:00011:00002",
  "USGS:11504115:00011:00010",
  "USGS:11504115:00011:00006",
  "USGS:11504115:00011:00003",
  "USGS:11504115:00011:00001",
  "USGS:11504115:00011:00009",
  "USGS:11504300:00011:00001",
  "USGS:11505800:00011:00001",
  "USGS:11505900:00011:00001",
  "USGS:11507000:00011:00001",
  "USGS:11507001:00011:00002",
  "USGS:412733081380500:00011:00007",
  "USGS:412733081380500:00011:00003",
  "USGS:412733081380500:00011:00004",
  "USGS:412733081380500:00011:00001",
  "USGS:412733081380500:00011:00005",
  "USGS:412733081380500:00011:00006",
  "USGS:412733081380500:00011:00008",
  "USGS:412743081381400:00011:00007",
  "USGS:412743081381400:00011:00003",
  "USGS:412743081381400:00011:00004",
  "USGS:412743081381400:00011:00001",
  "USGS:412743081381400:00011:00005",
  "USGS:412743081381400:00011:00008",
  "USGS:413108084415300:00011:00001",
  "USGS:414514081174400:00011:00006",
  "USGS:414514081174400:00011:00003",
  "USGS:414514081174400:00011:00004",
  "USGS:414514081174400:00011:00001",
  "USGS:414514081174400:00011:00009",
  "USGS:414514081174400:00011:00005",
  "USGS:414514081174400:00011:00007",
  "USGS:07185000:00011:00015",
  "USGS:07185000:00011:00005",
  "USGS:07185000:00011:00004",
  "USGS:07185080:00011:00014",
  "USGS:07185090:00011:00002",
  "USGS:07185090:00011:00001",
  "USGS:07185095:00011:00017",
  "USGS:07185095:00011:00001",
  "USGS:07185095:00011:00002",
  "USGS:07188000:00011:00015",
  "USGS:07188000:00011:00005",
  "USGS:07188000:00011:00016",
  "USGS:07189540:00011:00002",
  "USGS:07189540:00011:00001",
  "USGS:07189542:00011:00002",
  "USGS:07189542:00011:00001",
  "USGS:07190000:00011:00004",
  "USGS:07190000:00011:00003",
  "USGS:07190500:00011:00009",
  "USGS:07190500:00011:00008",
  "USGS:07191000:00011:00014",
  "USGS:07191000:00011:00004",
  "USGS:07191000:00011:00003",
  "USGS:07191220:00011:00005",
  "USGS:07191220:00011:00004",
  "USGS:07191220:00011:00003",
  "USGS:071912213:00011:00013",
  "USGS:01384500:00011:00001",
  "USGS:01384500:00011:00002",
  "USGS:01386000:00011:00001",
  "USGS:01386000:00011:00013",
  "USGS:01386990:00011:00001",
  "USGS:01386990:00011:00002",
  "USGS:01387000:00011:00002",
  "USGS:01387000:00011:00003",
  "USGS:01387500:00011:00001",
  "USGS:01387500:00011:00004",
  "USGS:01387905:00011:00002",
  "USGS:01387940:00011:00002",
  "USGS:01387940:00011:00001",
  "USGS:01387998:00011:00013",
  "USGS:01387998:00011:00012",
  "USGS:01388000:00011:00020",
  "USGS:01388000:00011:00001",
  "USGS:01388000:00011:00003",
  "USGS:01388000:00011:00021",
  "USGS:01388000:00011:00022",
  "USGS:01388000:00011:00033",
  "USGS:01388000:00011:00034",
  "USGS:01388100:00011:00002",
  "USGS:01388100:00011:00001",
  "USGS:01388500:00011:00001",
  "USGS:01388500:00011:00002",
  "USGS:01388700:00011:00001",
  "USGS:01388910:00011:00001",
  "USGS:01389005:00011:00022",
  "USGS:07161450:00011:00004",
  "USGS:01389005:00011:00025",
  "USGS:01389005:00011:00028",
  "USGS:01389005:00011:00009",
  "USGS:01389005:00011:00023",
  "USGS:01389005:00011:00026",
  "USGS:01389005:00011:00029",
  "USGS:01389005:00011:00024",
  "USGS:01389005:00011:00027",
  "USGS:01389005:00011:00030",
  "USGS:01389005:00011:00037",
  "USGS:01389005:00011:00038",
  "USGS:01389005:00011:00039",
  "USGS:01389005:00011:00040",
  "USGS:01389005:00011:00041",
  "USGS:01389005:00011:00042",
  "USGS:01389005:00011:00049",
  "USGS:01389005:00011:00050",
  "USGS:01389005:00011:00061",
  "USGS:01389005:00011:00062",
  "USGS:01389005:00011:00063",
  "USGS:01389005:00011:00043",
  "USGS:01389005:00011:00045",
  "USGS:01389010:00011:00002",
  "USGS:01389492:00011:00001",
  "USGS:01389500:00011:00002",
  "USGS:01389500:00011:00007",
  "USGS:01389534:00011:00001",
  "USGS:01389550:00011:00001",
  "USGS:01389550:00011:00002",
  "USGS:01389765:00011:00012",
  "USGS:01389765:00011:00001",
  "USGS:01389802:00011:00002",
  "USGS:01389890:00011:00002",
  "USGS:01389890:00011:00001",
  "USGS:01390450:00011:00013",
  "USGS:01390450:00011:00002",
  "USGS:01390450:00011:00001",
  "USGS:01390500:00011:00001",
  "USGS:01390500:00011:00002",
  "USGS:01391000:00011:00001",
  "USGS:01391000:00011:00002",
  "USGS:01391102:00011:00001",
  "USGS:01391102:00011:00002",
  "USGS:01391500:00011:00001",
  "USGS:01391500:00011:00002",
  "USGS:01392170:00011:00001",
  "USGS:01392500:00011:00001",
  "USGS:01392500:00011:00002",
  "USGS:01392650:00011:00005",
  "USGS:01392650:00011:00001",
  "USGS:01393450:00011:00001",
  "USGS:01393450:00011:00002",
  "USGS:01393890:00011:00004",
  "USGS:01393890:00011:00001",
  "USGS:01393895:00011:00002",
  "USGS:01393895:00011:00001",
  "USGS:01394000:00011:00002",
  "USGS:01394500:00011:00001",
  "USGS:01394500:00011:00002",
  "USGS:01394500:00011:00019",
  "USGS:01394620:00011:00011",
  "USGS:01394620:00011:00001",
  "USGS:01395000:00011:00001",
  "USGS:01395000:00011:00002",
  "USGS:01396000:00011:00002",
  "USGS:01396091:00011:00002",
  "USGS:01396091:00011:00001",
  "USGS:01396152:00011:00001",
  "USGS:01396152:00011:00002",
  "USGS:01396500:00011:00005",
  "USGS:01396500:00011:00007",
  "USGS:01396582:00011:00004",
  "USGS:01396582:00011:00001",
  "USGS:01396582:00011:00002",
  "USGS:01396660:00011:00001",
  "USGS:01396660:00011:00002",
  "USGS:01396790:00011:00002",
  "USGS:01396790:00011:00001",
  "USGS:01396800:00011:00002",
  "USGS:01396800:00011:00003",
  "USGS:01397000:00011:00002",
  "USGS:01397000:00011:00006",
  "USGS:01397420:00011:00001",
  "USGS:01398000:00011:00001",
  "USGS:01398000:00011:00002",
  "USGS:01398102:00011:00001",
  "USGS:02248600:00011:00003",
  "USGS:403541075112301:00011:00001",
  "USGS:403644074352701:00011:00001",
  "USGS:403719075091801:00011:00001",
  "USGS:403811074270501:00011:00001",
  "USGS:403824074545601:00011:00001",
  "USGS:404014074585401:00011:00001",
  "USGS:404059074223301:00011:00001",
  "USGS:404106074171901:00011:00001",
  "USGS:404217074294701:00011:00002",
  "USGS:404218074413701:00011:00001",
  "USGS:404223074381101:00011:00001",
  "USGS:404247074072301:00011:00002",
  "USGS:404405074161401:00011:00001",
  "USGS:404550074171600:00011:00001",
  "USGS:404751074250601:00011:00002",
  "USGS:404822074442601:00011:00001",
  "USGS:404934074400501:00011:00001",
  "USGS:404955074171101:00011:00002",
  "USGS:405002074310001:00011:00002",
  "USGS:405030074380901:00011:00002",
  "USGS:405219074132001:00011:00001",
  "USGS:405236074051801:00011:00002",
  "USGS:405305074105401:00011:00002",
  "USGS:405343074235201:00011:00002",
  "USGS:405424074355001:00011:00002",
  "USGS:405437074151001:00011:00002",
  "USGS:405502074395601:00011:00001",
  "USGS:405529074180901:00011:00002",
  "USGS:405658074332601:00011:00001",
  "USGS:405811074165501:00011:00002",
  "USGS:405934074120201:00011:00002",
  "USGS:405934074164401:00011:00001",
  "USGS:405939074084301:00011:00002",
  "USGS:410043074025301:00011:00001",
  "USGS:410139074150001:00011:00002",
  "USGS:410148074252901:00011:00002",
  "USGS:410207074270001:00011:00001",
  "USGS:410212074022101:00011:00001",
  "USGS:410230074300001:00011:00002",
  "USGS:410239074173501:00011:00002",
  "USGS:07324300:00011:00014",
  "USGS:07324300:00011:00004",
  "USGS:07324300:00011:00003",
  "USGS:07324400:00011:00007",
  "USGS:07324400:00011:00006",
  "USGS:07324400:00011:00005",
  "USGS:07325000:00011:00016",
  "USGS:07325000:00011:00006",
  "USGS:07325000:00011:00005",
  "USGS:07325500:00011:00018",
  "USGS:07325500:00011:00020",
  "USGS:07325500:00011:00019",
  "USGS:07325800:00011:00005",
  "USGS:07325800:00011:00004",
  "USGS:07325800:00011:00003",
  "USGS:07325840:00011:00003",
  "USGS:07325840:00011:00002",
  "USGS:07325840:00011:00001",
  "USGS:01429500:00011:00001",
  "USGS:01429500:00011:00002",
  "USGS:01430000:00011:00003",
  "USGS:01430000:00011:00001",
  "USGS:01430000:00011:00002",
  "USGS:01431500:00011:00017",
  "USGS:01431500:00011:00003",
  "USGS:01431500:00011:00001",
  "USGS:01431500:00011:00002",
  "USGS:01432110:00011:00012",
  "USGS:01432110:00011:00002",
  "USGS:01432110:00011:00001",
  "USGS:01432160:00011:00001",
  "USGS:01432160:00011:00003",
  "USGS:01432805:00011:00001",
  "USGS:01434000:00011:00005",
  "USGS:01434000:00011:00002",
  "USGS:01438500:00011:00004",
  "USGS:01438500:00011:00005",
  "USGS:01439500:00011:00004",
  "USGS:01439500:00011:00003",
  "USGS:01439590:00011:00002",
  "USGS:01439590:00011:00001",
  "USGS:01440400:00011:00004",
  "USGS:01440400:00011:00003",
  "USGS:01440485:00011:00002",
  "USGS:01440485:00011:00001",
  "USGS:01441495:00011:00002",
  "USGS:01441495:00011:00001",
  "USGS:07161450:00011:00014",
  "USGS:07161450:00011:00003",
  "USGS:07164500:00011:00014",
  "USGS:07164500:00011:00012",
  "USGS:07164500:00011:00011",
  "USGS:07164500:00011:00030",
  "USGS:07164600:00011:00004",
  "USGS:07164600:00011:00003",
  "USGS:07165562:00011:00004",
  "USGS:07165562:00011:00003",
  "USGS:07165565:00011:00004",
  "USGS:07165565:00011:00003",
  "USGS:07165570:00011:00005",
  "USGS:07165570:00011:00004",
  "USGS:07165570:00011:00003",
  "USGS:07171000:00011:00006",
  "USGS:07171000:00011:00005",
  "USGS:07174400:00011:00014",
  "USGS:07174400:00011:00004",
  "USGS:07174400:00011:00003",
  "USGS:07174470:00011:00014",
  "USGS:07174470:00011:00002",
  "USGS:07174470:00011:00001",
  "USGS:07174618:00011:00003",
  "USGS:07174618:00011:00001",
  "USGS:07175500:00011:00016",
  "USGS:07175500:00011:00006",
  "USGS:07175500:00011:00005",
  "USGS:07176000:00011:00005",
  "USGS:07176000:00011:00004",
  "USGS:07176321:00011:00005",
  "USGS:07176500:00011:00014",
  "USGS:07176500:00011:00004",
  "USGS:07176500:00011:00003",
  "USGS:07176950:00011:00014",
  "USGS:07176950:00011:00002",
  "USGS:07176950:00011:00001",
  "USGS:07177500:00011:00019",
  "USGS:07177500:00011:00018",
  "USGS:07177500:00011:00008",
  "USGS:07177500:00011:00007",
  "USGS:07177500:00011:00020",
  "USGS:07177500:00011:00022",
  "USGS:07177500:00011:00021",
  "USGS:07177650:00011:00004",
  "USGS:07177650:00011:00003",
  "USGS:07177800:00011:00004",
  "USGS:07177800:00011:00003",
  "USGS:07178000:00011:00008",
  "USGS:07178000:00011:00007",
  "USGS:07178200:00011:00009",
  "USGS:07178200:00011:00008",
  "USGS:07178200:00011:00007",
  "USGS:07178200:00011:00010",
  "USGS:07178200:00011:00012",
  "USGS:07178200:00011:00011",
  "USGS:07178452:00011:00003",
  "USGS:07178452:00011:00001",
  "USGS:07178645:00011:00003",
  "USGS:07178645:00011:00001",
  "USGS:410449074483301:00011:00001",
  "USGS:410622074570901:00011:00001",
  "USGS:410639074293001:00011:00002",
  "USGS:410716074141601:00011:00002",
  "USGS:410800074204301:00011:00002",
  "USGS:410811074182801:00011:00002",
  "USGS:410914074540401:00011:00001",
  "USGS:410946074403101:00011:00001",
  "USGS:411130074252501:00011:00002",
  "USGS:01109403:00011:00002",
  "USGS:01109403:00011:00001",
  "USGS:01111300:00011:00001",
  "USGS:01111300:00011:00002",
  "USGS:01111500:00011:00001",
  "USGS:01111500:00011:00002",
  "USGS:01112500:00011:00002",
  "USGS:01112500:00011:00016",
  "USGS:01113895:00011:00001",
  "USGS:01113895:00011:00002",
  "USGS:01114000:00011:00001",
  "USGS:01114000:00011:00003",
  "USGS:01114500:00011:00001",
  "USGS:01114500:00011:00003",
  "USGS:01115098:00011:00004",
  "USGS:01115098:00011:00003",
  "USGS:01115098:00011:00001",
  "USGS:01115098:00011:00002",
  "USGS:01115110:00011:00002",
  "USGS:01115110:00011:00004",
  "USGS:01115110:00011:00001",
  "USGS:071912213:00011:00003",
  "USGS:071912213:00011:00002",
  "USGS:071912213:00011:00001",
  "USGS:071912213:00011:00014",
  "USGS:071912213:00011:00016",
  "USGS:071912213:00011:00015",
  "USGS:071912213:00011:00017",
  "USGS:07191222:00011:00014",
  "USGS:07191222:00011:00002",
  "USGS:07191222:00011:00001",
  "USGS:07191222:00011:00015",
  "USGS:07191222:00011:00016",
  "USGS:07191222:00011:00017",
  "USGS:07191222:00011:00018",
  "USGS:07191285:00011:00003",
  "USGS:07191285:00011:00002",
  "USGS:07191285:00011:00001",
  "USGS:07191288:00011:00003",
  "USGS:07191288:00011:00002",
  "USGS:07191288:00011:00001",
  "USGS:07191300:00011:00016",
  "USGS:07191300:00011:00004",
  "USGS:07191300:00011:00003",
  "USGS:07191400:00011:00015",
  "USGS:07191400:00011:00004",
  "USGS:07191400:00011:00003",
  "USGS:07191500:00011:00005",
  "USGS:07191500:00011:00004",
  "USGS:07194500:00011:00003",
  "USGS:07194500:00011:00017",
  "USGS:07194500:00011:00016",
  "USGS:07194555:00011:00003",
  "USGS:07194555:00011:00001",
  "USGS:07195500:00011:00014",
  "USGS:07195500:00011:00004",
  "USGS:07195500:00011:00003",
  "USGS:07195855:00011:00013",
  "USGS:07195855:00011:00002",
  "USGS:07195855:00011:00001",
  "USGS:07195865:00011:00002",
  "USGS:07195865:00011:00001",
  "USGS:07196000:00011:00014",
  "USGS:07196000:00011:00004",
  "USGS:07196000:00011:00003",
  "USGS:07196090:00011:00004",
  "USGS:07196090:00011:00002",
  "USGS:07196090:00011:00001",
  "USGS:07196500:00011:00014",
  "USGS:07196500:00011:00004",
  "USGS:07196500:00011:00003",
  "USGS:07197000:00011:00014",
  "USGS:07197000:00011:00004",
  "USGS:07197000:00011:00015",
  "USGS:07197360:00011:00018",
  "USGS:07197360:00011:00002",
  "USGS:07197360:00011:00016",
  "USGS:07198000:00011:00001",
  "USGS:07198000:00011:00016",
  "USGS:07198000:00011:00019",
  "USGS:07198000:00011:00018",
  "USGS:07198000:00011:00021",
  "USGS:07228500:00011:00008",
  "USGS:07228500:00011:00019",
  "USGS:07228940:00011:00002",
  "USGS:07228940:00011:00001",
  "USGS:07229050:00011:00002",
  "USGS:07229050:00011:00015",
  "USGS:07229200:00011:00016",
  "USGS:07229200:00011:00006",
  "USGS:07229200:00011:00005",
  "USGS:07229445:00011:00015",
  "USGS:07229445:00011:00002",
  "USGS:07229445:00011:00001",
  "USGS:07229445:00011:00014",
  "USGS:07229900:00011:00005",
  "USGS:07229900:00011:00004",
  "USGS:07230000:00011:00007",
  "USGS:07230000:00011:00006",
  "USGS:07230500:00011:00004",
  "USGS:07230500:00011:00003",
  "USGS:07231000:00011:00007",
  "USGS:07231000:00011:00006",
  "USGS:07231500:00011:00016",
  "USGS:07231500:00011:00006",
  "USGS:07231500:00011:00017",
  "USGS:07232470:00011:00003",
  "USGS:07232470:00011:00014",
  "USGS:07232470:00011:00013",
  "USGS:07234000:00011:00016",
  "USGS:07234000:00011:00006",
  "USGS:07234000:00011:00005",
  "USGS:07235600:00011:00003",
  "USGS:07235600:00011:00002",
  "USGS:07235600:00011:00001",
  "USGS:07237500:00011:00017",
  "USGS:07237500:00011:00006",
  "USGS:07237500:00011:00005",
  "USGS:07238000:00011:00014",
  "USGS:07238000:00011:00004",
  "USGS:07238000:00011:00003",
  "USGS:07238500:00011:00022",
  "USGS:07238500:00011:00021",
  "USGS:07239000:00011:00017",
  "USGS:07239000:00011:00016",
  "USGS:07239300:00011:00014",
  "USGS:07239300:00011:00004",
  "USGS:07239300:00011:00003",
  "USGS:07239450:00011:00009",
  "USGS:07239450:00011:00008",
  "USGS:07239450:00011:00007",
  "USGS:07239450:00011:00010",
  "USGS:07239450:00011:00021",
  "USGS:07239450:00011:00011",
  "USGS:07239500:00011:00026",
  "USGS:07239500:00011:00016",
  "USGS:07239500:00011:00006",
  "USGS:07239500:00011:00005",
  "USGS:07239500:00011:00027",
  "USGS:07239700:00011:00001",
  "USGS:07239700:00011:00005",
  "USGS:07239700:00011:00004",
  "USGS:07239700:00011:00006",
  "USGS:01115190:00011:00002",
  "USGS:01115110:00011:00003",
  "USGS:01115114:00011:00003",
  "USGS:01115114:00011:00002",
  "USGS:01115114:00011:00001",
  "USGS:01115114:00011:00004",
  "USGS:01115120:00011:00003",
  "USGS:01115120:00011:00002",
  "USGS:01115120:00011:00001",
  "USGS:01115120:00011:00004",
  "USGS:01115170:00011:00002",
  "USGS:01115170:00011:00004",
  "USGS:01115170:00011:00001",
  "USGS:01115170:00011:00003",
  "USGS:01115183:00011:00002",
  "USGS:01115183:00011:00004",
  "USGS:01115183:00011:00001",
  "USGS:01115183:00011:00003",
  "USGS:01115184:00011:00003",
  "USGS:01115184:00011:00002",
  "USGS:01115184:00011:00001",
  "USGS:01115184:00011:00004",
  "USGS:01115187:00011:00015",
  "USGS:01115187:00011:00017",
  "USGS:01115187:00011:00016",
  "USGS:01115187:00011:00003",
  "USGS:01115187:00011:00002",
  "USGS:01115187:00011:00014",
  "USGS:0208111310:00011:00002",
  "USGS:0208111310:00011:00001",
  "USGS:340643095044801:00011:00001",
  "USGS:340643095044801:00011:00002",
  "USGS:340643095044801:00011:00003",
  "USGS:340643095044801:00011:00004",
  "USGS:340643095044801:00011:00005",
  "USGS:340643095044801:00011:00006",
  "USGS:340643095044801:00011:00007",
  "USGS:342527096493301:00011:00001",
  "USGS:342633096494401:00011:00001",
  "USGS:343017096561501:00011:00002",
  "USGS:343017096561501:00011:00001",
  "USGS:343022096565701:00011:00001",
  "USGS:343457096404501:00011:00001",
  "USGS:344749098350301:00011:00001",
  "USGS:345759099163401:00011:00001",
  "USGS:350748098231101:00011:00001",
  "USGS:350755099283201:00011:00001",
  "USGS:351223099480001:00011:00001",
  "USGS:351308098341601:00011:00001",
  "USGS:351521099522901:00011:00001",
  "USGS:351727098290401:00011:00001",
  "USGS:352423098341701:00011:00001",
  "USGS:352523097032101:00011:00002",
  "USGS:352523097032101:00011:00003",
  "USGS:352523097032101:00011:00001",
  "USGS:352537099234301:00011:00011",
  "USGS:352537099234301:00011:00001",
  "USGS:352802098191601:00011:00001",
  "USGS:352959097114001:00011:00002",
  "USGS:352959097114001:00011:00001",
  "USGS:353002097114001:00011:00002",
  "USGS:353002097114001:00011:00001",
  "USGS:353211098191501:00011:00002",
  "USGS:353211098191501:00011:00001",
  "USGS:355133099434901:00011:00001",
  "USGS:355510096293501:00011:00001",
  "USGS:361739099323301:00011:00001",
  "USGS:362823096224201:00011:00001",
  "USGS:363021096432402:00011:00001",
  "USGS:363021096432403:00011:00003",
  "USGS:363021096432403:00011:00001",
  "USGS:363021096432404:00011:00001",
  "USGS:363033101440701:00011:00001",
  "USGS:364001096184901:00011:00001",
  "USGS:364001096184903:00011:00001",
  "USGS:364821098144901:00011:00001",
  "USGS:364831098120201:00011:00002",
  "USGS:364831098120201:00011:00001",
  "USGS:365942094504203:00011:00001",
  "USGS:0208758850:00011:00002",
  "USGS:0208758850:00011:00001",
  "USGS:0208773375:00011:00011",
  "USGS:0208773375:00011:00001",
  "USGS:02088000:00011:00001",
  "USGS:02088000:00011:00002",
  "USGS:02088383:00011:00002",
  "USGS:02088383:00011:00001",
  "USGS:394808075172401:00011:00001",
  "USGS:394808075172402:00011:00001",
  "USGS:394808075172404:00011:00001",
  "USGS:394829074053503:00011:00001",
  "USGS:394957075053001:00011:00001",
  "USGS:395150074284201:00011:00001",
  "USGS:395206075111801:00011:   NA",
  "USGS:395315074494601:00011:00001",
  "USGS:395343074492501:00011:00001",
  "USGS:395524074502501:00011:00001",
  "USGS:395524074502502:00011:00001",
  "USGS:395525074502505:00011:00001",
  "USGS:395525074502601:00011:00001",
  "USGS:395609074124001:00011:00001",
  "USGS:395722074374001:00011:00001",
  "USGS:395928074502701:00011:00001",
  "USGS:395930074142101:00011:00001",
  "USGS:400210074031001:00011:00001",
  "USGS:400210074031002:00011:00001",
  "USGS:400232074213201:00011:00001",
  "USGS:400530074090901:00011:00001",
  "USGS:400642074024101:00011:00003",
  "USGS:400642074024101:00011:00005",
  "USGS:400642074024101:00011:00006",
  "USGS:400642074024101:00011:00008",
  "USGS:400642074024101:00011:00002",
  "USGS:400642074024101:00011:00004",
  "USGS:400642074024101:00011:00007",
  "USGS:400711074020201:00011:00001",
  "USGS:400832074082101:00011:00001",
  "USGS:401105074120201:00011:00001",
  "USGS:401105074120202:00011:00001",
  "USGS:401105074120204:00011:00001",
  "USGS:401105074120205:00011:00001",
  "USGS:401542074053001:00011:00001",
  "USGS:401552074501801:00011:00001",
  "USGS:401616074462401:00011:00001",
  "USGS:401804074432601:00011:00001",
  "USGS:401834074515501:00011:00001",
  "USGS:402109074301301:00011:00001",
  "USGS:402109074301302:00011:00001",
  "USGS:402138074435801:00011:00001",
  "USGS:402143074185201:00011:00001",
  "USGS:402151074525301:00011:00001",
  "USGS:402414074584401:00011:00001",
  "USGS:402454074205601:00011:00001",
  "USGS:402504074414201:00011:00001",
  "USGS:402512074414301:00011:00001",
  "USGS:402553074271701:00011:00001",
  "USGS:402644074563601:00011:00001",
  "USGS:402657074085101:00011:00002",
  "USGS:402657074085101:00011:00004",
  "USGS:402657074085101:00011:00005",
  "USGS:402657074085101:00011:00007",
  "USGS:402657074085101:00011:00001",
  "USGS:402657074085101:00011:00003",
  "USGS:402657074085101:00011:00006",
  "USGS:402758074431301:00011:00001",
  "USGS:02102500:00011:00004",
  "USGS:02102500:00011:00005",
  "USGS:02102908:00011:00001",
  "USGS:02102908:00011:00002",
  "USGS:02102908:00011:00003",
  "USGS:02103000:00011:00001",
  "USGS:02103000:00011:00002",
  "USGS:02104000:00011:00002",
  "USGS:02104220:00011:00002",
  "USGS:02104220:00011:00001",
  "USGS:02105500:00011:00016",
  "USGS:02105500:00011:00002",
  "USGS:02105500:00011:00003",
  "USGS:02105769:00011:   NA",
  "USGS:02105769:00011:   NA",
  "USGS:02105769:00011:   NA",
  "USGS:02106500:00011:00002",
  "USGS:02106500:00011:00003",
  "USGS:02108000:00011:00002",
  "USGS:02108000:00011:00003",
  "USGS:02108566:00011:00003",
  "USGS:02109500:00011:00002",
  "USGS:02109500:00011:00003",
  "USGS:02111000:00011:00016",
  "USGS:02111000:00011:00005",
  "USGS:02111000:00011:00001",
  "USGS:02111000:00011:00002",
  "USGS:02111180:00011:00005",
  "USGS:02111180:00011:00001",
  "USGS:02111180:00011:00002",
  "USGS:02111391:00011:00002",
  "USGS:01463620:00011:00002",
  "USGS:01463740:00011:00002",
  "USGS:01463740:00011:00001",
  "USGS:01463882:00011:00001",
  "USGS:01464000:00011:00001",
  "USGS:01464000:00011:00002",
  "USGS:01464500:00011:00002",
  "USGS:01464500:00011:00005",
  "USGS:01465850:00011:00004",
  "USGS:01465850:00011:00003",
  "USGS:01465880:00011:00001",
  "USGS:01466500:00011:00001",
  "USGS:01466500:00011:00002",
  "USGS:01466500:00011:00006",
  "USGS:01466900:00011:00020",
  "USGS:01466900:00011:00002",
  "USGS:01466900:00011:00001",
  "USGS:01467000:00011:00001",
  "USGS:01467000:00011:00002",
  "USGS:01467005:00011:00001",
  "USGS:01467081:00011:00001",
  "USGS:01467081:00011:00002",
  "USGS:01467150:00011:00002",
  "USGS:01467150:00011:00018",
  "USGS:01475001:00011:00002",
  "USGS:01475001:00011:00001",
  "USGS:01477120:00011:00018",
  "USGS:01477120:00011:00002",
  "USGS:01477120:00011:00005",
  "USGS:01482500:00011:00001",
  "USGS:01482500:00011:00002",
  "USGS:04253400:00011:00002",
  "USGS:385655074532601:00011:00002",
  "USGS:385655074532601:00011:00004",
  "USGS:385655074532601:00011:00005",
  "USGS:385655074532601:00011:00007",
  "USGS:385655074532601:00011:00001",
  "USGS:385655074532601:00011:00003",
  "USGS:385655074532601:00011:00006",
  "USGS:385709074512801:00011:00001",
  "USGS:385804074574201:00011:00001",
  "USGS:390002074541002:00011:00001",
  "USGS:390012074472001:00011:00001",
  "USGS:390156074533401:00011:00001",
  "USGS:390422074544701:00011:00001",
  "USGS:390425074544601:00011:00001",
  "USGS:390608074483801:00011:00001",
  "USGS:391827074371001:00011:00001",
  "USGS:392017074300201:00011:00001",
  "USGS:392032074300801:00011:00001",
  "USGS:392239074252401:00011:00002",
  "USGS:392239074252401:00011:00004",
  "USGS:392239074252401:00011:00005",
  "USGS:392239074252401:00011:00007",
  "USGS:392239074252401:00011:00001",
  "USGS:392239074252401:00011:00003",
  "USGS:392239074252401:00011:00006",
  "USGS:392245075211901:00011:00001",
  "USGS:392731075092401:00011:00001",
  "USGS:392732075092401:00011:00001",
  "USGS:392754074270101:00011:00001",
  "USGS:393232074263901:00011:00001",
  "USGS:393232074263903:00011:00001",
  "USGS:393333074442401:00011:00001",
  "USGS:393348075275701:00011:00001",
  "USGS:393541074510601:00011:00001",
  "USGS:393838075194901:00011:00001",
  "USGS:394037075191501:00011:00001",
  "USGS:394119075062701:00011:00001",
  "USGS:394215074561701:00011:00001",
  "USGS:394215074561702:00011:00001",
  "USGS:394215074561703:00011:00001",
  "USGS:394221075072201:00011:00001",
  "USGS:394236075272101:00011:00001",
  "USGS:394256075101001:00011:00001",
  "USGS:394354075025901:00011:00001",
  "USGS:394540074062901:00011:00002",
  "USGS:394540074062901:00011:00004",
  "USGS:394540074062901:00011:00005",
  "USGS:394540074062901:00011:00007",
  "USGS:394540074062901:00011:00001",
  "USGS:394540074062901:00011:00006",
  "USGS:02146750:00011:00006",
  "USGS:02146750:00011:00001",
  "USGS:02146750:00011:00002",
  "USGS:0214678175:00011:00002",
  "USGS:01411300:00011:00002",
  "USGS:01411300:00011:00003",
  "USGS:01411320:00011:00005",
  "USGS:01411320:00011:00001",
  "USGS:01411330:00011:00005",
  "USGS:01411330:00011:00001",
  "USGS:01411350:00011:00015",
  "USGS:01411350:00011:00001",
  "USGS:01411355:00011:00015",
  "USGS:01411355:00011:00001",
  "USGS:01411360:00011:00015",
  "USGS:01411360:00011:00001",
  "USGS:01411390:00011:00004",
  "USGS:01411390:00011:00001",
  "USGS:01411435:00011:00015",
  "USGS:01411435:00011:00001",
  "USGS:01411456:00011:00002",
  "USGS:01411456:00011:00001",
  "USGS:01411500:00011:00002",
  "USGS:01411500:00011:00006",
  "USGS:01412150:00011:00001",
  "USGS:01412800:00011:00001",
  "USGS:01412800:00011:00002",
  "USGS:01413038:00011:00015",
  "USGS:01413038:00011:00002",
  "USGS:01439800:00011:00001",
  "USGS:01439800:00011:00002",
  "USGS:01440000:00011:00001",
  "USGS:01440000:00011:00002",
  "USGS:01440200:00011:00019",
  "USGS:01440200:00011:00002",
  "USGS:01443280:00011:00002",
  "USGS:01443280:00011:00001",
  "USGS:01443500:00011:00001",
  "USGS:01443500:00011:00002",
  "USGS:01443900:00011:00001",
  "USGS:01443900:00011:00002",
  "USGS:01445000:00011:00001",
  "USGS:01445000:00011:00002",
  "USGS:01445500:00011:00001",
  "USGS:01445500:00011:00002",
  "USGS:01446000:00011:00001",
  "USGS:01446000:00011:00002",
  "USGS:01446500:00011:00001",
  "USGS:01446500:00011:00002",
  "USGS:01446995:00011:00001",
  "USGS:01455090:00011:00002",
  "USGS:01455090:00011:00001",
  "USGS:01455400:00011:00002",
  "USGS:01455400:00011:00001",
  "USGS:01455500:00011:00001",
  "USGS:01455500:00011:00002",
  "USGS:01457000:00011:00001",
  "USGS:01457000:00011:00002",
  "USGS:01457500:00011:00003",
  "USGS:01458500:00011:00013",
  "USGS:01458500:00011:00001",
  "USGS:01458500:00011:00015",
  "USGS:01458500:00011:00017",
  "USGS:01458500:00011:00016",
  "USGS:01458500:00011:00014",
  "USGS:01458500:00011:00018",
  "USGS:01460440:00011:00003",
  "USGS:01460440:00011:00011",
  "USGS:01460440:00011:00009",
  "USGS:01460595:00011:00002",
  "USGS:01460595:00011:00003",
  "USGS:01460595:00011:00004",
  "USGS:01460595:00011:00005",
  "USGS:01460880:00011:00002",
  "USGS:01460880:00011:00003",
  "USGS:01461500:00011:00001",
  "USGS:01462000:00011:00015",
  "USGS:01462000:00011:00002",
  "USGS:01462500:00011:00001",
  "USGS:01463500:00011:00009",
  "USGS:01463500:00011:00005",
  "USGS:01463500:00011:00012",
  "USGS:01463500:00011:00026",
  "USGS:01463500:00011:00028",
  "USGS:01463500:00011:00027",
  "USGS:01463500:00011:00025",
  "USGS:01463500:00011:00031",
  "USGS:02137727:00011:00018",
  "USGS:02137727:00011:00016",
  "USGS:02137727:00011:00001",
  "USGS:02137727:00011:00002",
  "USGS:02138500:00011:00001",
  "USGS:02138500:00011:00002",
  "USGS:02138520:00011:00011",
  "USGS:02248600:00011:00001",
  "USGS:02248600:00011:00005",
  "USGS:02248600:00011:00004",
  "USGS:07240000:00011:00004",
  "USGS:07240000:00011:00003",
  "USGS:07240200:00011:00001",
  "USGS:07240500:00011:00005",
  "USGS:07240500:00011:00004",
  "USGS:07241000:00011:00015",
  "USGS:07241000:00011:00031",
  "USGS:07241000:00011:00004",
  "USGS:07241000:00011:00003",
  "USGS:07241000:00011:00014",
  "USGS:07241000:00011:00017",
  "USGS:07241000:00011:00008",
  "USGS:07241520:00011:00004",
  "USGS:07241520:00011:00002",
  "USGS:07241520:00011:00023",
  "USGS:07241520:00011:00003",
  "USGS:07241520:00011:00006",
  "USGS:07241550:00011:00018",
  "USGS:07241550:00011:00006",
  "USGS:07241550:00011:00012",
  "USGS:07241550:00011:00019",
  "USGS:07241550:00011:00021",
  "USGS:07241550:00011:00020",
  "USGS:07241588:00011:00003",
  "USGS:07241588:00011:00001",
  "USGS:07241600:00011:00002",
  "USGS:07241600:00011:00014",
  "USGS:07241600:00011:00015",
  "USGS:07241600:00011:00019",
  "USGS:07241600:00011:00001",
  "USGS:07241600:00011:00013",
  "USGS:07241600:00011:00017",
  "USGS:07241600:00011:00016",
  "USGS:07241800:00011:00002",
  "USGS:07241800:00011:00001",
  "USGS:07242000:00011:00017",
  "USGS:07242000:00011:00007",
  "USGS:07242000:00011:00018",
  "USGS:07242380:00011:00004",
  "USGS:07242380:00011:00003",
  "USGS:07243500:00011:00016",
  "USGS:07243500:00011:00006",
  "USGS:07243500:00011:00005",
  "USGS:07245000:00011:00023",
  "USGS:07245000:00011:00013",
  "USGS:07245000:00011:00012",
  "USGS:07246500:00011:00006",
  "USGS:07246500:00011:00004",
  "USGS:07247015:00011:00004",
  "USGS:07247015:00011:00003",
  "USGS:07247250:00011:00003",
  "USGS:07247250:00011:00002",
  "USGS:07247250:00011:00001",
  "USGS:07247500:00011:00005",
  "USGS:07247500:00011:00004",
  "USGS:07247500:00011:00003",
  "USGS:07249413:00011:00003",
  "USGS:07249413:00011:00002",
  "USGS:07249413:00011:00001",
  "USGS:07249800:00011:00022",
  "USGS:07249800:00011:00002",
  "USGS:07249800:00011:00001",
  "USGS:07249920:00011:00004",
  "USGS:07249920:00011:00001",
  "USGS:07249985:00011:00012",
  "USGS:07249985:00011:00011",
  "USGS:07249985:00011:00001",
  "USGS:07300500:00011:00006",
  "USGS:07300500:00011:00005",
  "USGS:07300500:00011:00004",
  "USGS:07301110:00011:00006",
  "USGS:07301110:00011:00005",
  "USGS:07301420:00011:00005",
  "USGS:07301420:00011:00004",
  "USGS:07301420:00011:00003",
  "USGS:07301481:00011:00014",
  "USGS:07301481:00011:00015",
  "USGS:07301500:00011:00001",
  "USGS:07301500:00011:00025",
  "USGS:07301500:00011:00015",
  "USGS:07301500:00011:00014",
  "USGS:07301500:00011:00003",
  "USGS:07302500:00011:00015",
  "USGS:07302500:00011:00004",
  "USGS:07302500:00011:00003",
  "USGS:07303000:00011:00004",
  "USGS:07303000:00011:00003",
  "USGS:07303400:00011:00001",
  "USGS:07303400:00011:00014",
  "USGS:07303400:00011:00013",
  "USGS:07303400:00011:00012",
  "USGS:07303400:00011:00003",
  "USGS:07303400:00011:00018",
  "USGS:07305000:00011:00001",
  "USGS:07305000:00011:00014",
  "USGS:07305000:00011:00013",
  "USGS:07305000:00011:00012",
  "USGS:07305000:00011:00003",
  "USGS:07307010:00011:00014",
  "USGS:07307010:00011:00016",
  "USGS:07307010:00011:00015",
  "USGS:07307028:00011:00016",
  "USGS:07307028:00011:00015",
  "USGS:07308990:00011:00002",
  "USGS:07308990:00011:00001",
  "USGS:07309435:00011:00013",
  "USGS:07309435:00011:00002",
  "USGS:07309435:00011:00001",
  "USGS:07309500:00011:00002",
  "USGS:07309500:00011:00001",
  "USGS:07309990:00011:00001",
  "USGS:07309990:00011:00003",
  "USGS:07311000:00011:00007",
  "USGS:07311000:00011:00006",
  "USGS:07311000:00011:00005",
  "USGS:07311230:00011:00001",
  "USGS:07311230:00011:00003",
  "USGS:07311240:00011:00001",
  "USGS:07311240:00011:00003",
  "USGS:07311415:00011:00003",
  "USGS:07311415:00011:00002",
  "USGS:07311415:00011:00001",
  "USGS:07311500:00011:00007",
  "USGS:07311500:00011:00006",
  "USGS:07312920:00011:00003",
  "USGS:07312920:00011:00001",
  "USGS:07313000:00011:00005",
  "USGS:07313000:00011:00003",
  "USGS:07313585:00011:00003",
  "USGS:07313585:00011:00001",
  "USGS:07315500:00011:00003",
  "USGS:07315500:00011:00017",
  "USGS:07315500:00011:00001",
  "USGS:07315500:00011:00002",
  "USGS:07315700:00011:00015",
  "USGS:07315700:00011:00014",
  "USGS:07316000:00011:00016",
  "USGS:07316000:00011:00006",
  "USGS:07316000:00011:00025",
  "USGS:07316500:00011:00014",
  "USGS:07316500:00011:00004",
  "USGS:07316500:00011:00003",
  "USGS:07324200:00011:00015",
  "USGS:07324200:00011:00014",
  "USGS:07324200:00011:00013",
  "USGS:335631078003604:00011:00001",
  "USGS:335631078003605:00011:00001",
  "USGS:335631078003606:00011:00001",
  "USGS:335849078054301:00011:00001",
  "USGS:344520079281001:00011:00001",
  "USGS:07325850:00011:00005",
  "USGS:07325850:00011:00004",
  "USGS:07325850:00011:00003",
  "USGS:07325860:00011:00005",
  "USGS:07325860:00011:00004",
  "USGS:07325860:00011:00003",
  "USGS:07325900:00011:00014",
  "USGS:07325900:00011:00003",
  "USGS:07326000:00011:00006",
  "USGS:07326000:00011:00005",
  "USGS:07326500:00011:00016",
  "USGS:07326500:00011:00006",
  "USGS:07326500:00011:00005",
  "USGS:07327442:00011:00004",
  "USGS:07327442:00011:00003",
  "USGS:07327447:00011:00004",
  "USGS:07327447:00011:00003",
  "USGS:07327447:00011:00017",
  "USGS:07327550:00011:00004",
  "USGS:07327550:00011:00003",
  "USGS:07328100:00011:00019",
  "USGS:07328100:00011:00009",
  "USGS:07328100:00011:00020",
  "USGS:07328180:00011:00002",
  "USGS:07328180:00011:00001",
  "USGS:07328500:00011:00014",
  "USGS:07328500:00011:00004",
  "USGS:07328500:00011:00003",
  "USGS:07329605:00011:00004",
  "USGS:07329605:00011:00002",
  "USGS:07329605:00011:00001",
  "USGS:07329605:00011:00005",
  "USGS:07329610:00011:00013",
  "USGS:07329610:00011:00002",
  "USGS:07329610:00011:00001",
  "USGS:07329700:00011:00017",
  "USGS:07329780:00011:00003",
  "USGS:07329780:00011:00002",
  "USGS:07329780:00011:00001",
  "USGS:07329849:00011:00001",
  "USGS:07329849:00011:00002",
  "USGS:073298507:00011:00003",
  "USGS:073298507:00011:00004",
  "USGS:073298507:00011:00014",
  "USGS:07329852:00011:00002",
  "USGS:07329852:00011:00001",
  "USGS:07331000:00011:00001",
  "USGS:07331000:00011:00017",
  "USGS:07331000:00011:00007",
  "USGS:07331000:00011:00018",
  "USGS:07331000:00011:00003",
  "USGS:07331200:00011:00003",
  "USGS:07331200:00011:00002",
  "USGS:07331200:00011:00001",
  "USGS:07331295:00011:00001",
  "USGS:07331300:00011:00012",
  "USGS:07331300:00011:00002",
  "USGS:07331300:00011:00001",
  "USGS:07331383:00011:00003",
  "USGS:07331383:00011:00001",
  "USGS:07332390:00011:00015",
  "USGS:07332390:00011:00003",
  "USGS:07332390:00011:00002",
  "USGS:07332500:00011:00015",
  "USGS:07332500:00011:00005",
  "USGS:07332500:00011:00004",
  "USGS:07333010:00011:00015",
  "USGS:07333010:00011:00002",
  "USGS:07333010:00011:00001",
  "USGS:07333010:00011:00014",
  "USGS:07333900:00011:00002",
  "USGS:07333900:00011:00015",
  "USGS:07333900:00011:00014",
  "USGS:07333900:00011:00001",
  "USGS:07334000:00011:00015",
  "USGS:07334000:00011:00005",
  "USGS:07334000:00011:00004",
  "USGS:07334200:00011:00021",
  "USGS:07334200:00011:00004",
  "USGS:07334200:00011:00006",
  "USGS:07334200:00011:00003",
  "USGS:07334238:00011:00001",
  "USGS:07334238:00011:00003",
  "USGS:07334800:00011:00001",
  "USGS:07335300:00011:00006",
  "USGS:07335300:00011:00005",
  "USGS:07335300:00011:00004",
  "USGS:07335500:00011:00014",
  "USGS:07335500:00011:00004",
  "USGS:07335500:00011:00003",
  "USGS:07335700:00011:00016",
  "USGS:07335700:00011:00005",
  "USGS:07335700:00011:00004",
  "USGS:07335700:00011:00003",
  "USGS:07335775:00011:00017",
  "USGS:07335775:00011:00016",
  "USGS:07335790:00011:00014",
  "USGS:07335790:00011:00004",
  "USGS:07335790:00011:00003",
  "USGS:07336200:00011:00014",
  "USGS:07336200:00011:00004",
  "USGS:07336200:00011:00003",
  "USGS:07337300:00011:00003",
  "USGS:07337300:00011:00015",
  "USGS:07337900:00011:00014",
  "USGS:07337900:00011:00004",
  "USGS:07337900:00011:00003",
  "USGS:07338500:00011:00015",
  "USGS:07338500:00011:00005",
  "USGS:07338500:00011:00004",
  "USGS:07338750:00011:00005",
  "USGS:07338750:00011:00004",
  "USGS:07338750:00011:00003",
  "USGS:07339000:00011:00001",
  "USGS:07339000:00011:00017",
  "USGS:07339000:00011:00006",
  "USGS:07339000:00011:00005",
  "USGS:340042095051801:00011:00001",
  "USGS:340643095044601:00011:00001",
  "USGS:340643095044601:00011:00002",
  "USGS:340643095044601:00011:00003",
  "USGS:340643095044601:00011:00004",
  "USGS:340643095044601:00011:00005",
  "USGS:340643095044601:00011:00006",
  "USGS:340643095044601:00011:00007",
  "USGS:340643095044601:00011:00008",
  "USGS:340643095044601:00011:00009",
  "USGS:340643095044601:00011:00010",
  "USGS:340643095044601:00011:00011",
  "USGS:01115630:00011:00001",
  "USGS:01115630:00011:00002",
  "USGS:02110400:00011:00001",
  "USGS:02110400:00011:00012",
  "USGS:02110400:00011:00008",
  "USGS:02110400:00011:00010",
  "USGS:02110400:00011:00018",
  "USGS:02110400:00011:00002",
  "USGS:02110400:00011:00003",
  "USGS:02110400:00011:00004",
  "USGS:02110400:00011:00006",
  "USGS:02110500:00011:00017",
  "USGS:02110500:00011:00001",
  "USGS:02110500:00011:00002",
  "USGS:02110500:00011:00022",
  "USGS:02110500:00011:00018",
  "USGS:02110500:00011:00019",
  "USGS:02110500:00011:00021",
  "USGS:02110550:00011:00006",
  "USGS:02110550:00011:00013",
  "USGS:02110550:00011:00003",
  "USGS:04188433:00011:00001",
  "USGS:04188496:00011:00021",
  "USGS:04188496:00011:00003",
  "USGS:04188496:00011:00002",
  "USGS:04188496:00011:00001",
  "USGS:04188496:00011:00019",
  "USGS:04188496:00011:00020",
  "USGS:04188496:00011:00022",
  "USGS:04188496:00011:00023",
  "USGS:04188496:00011:00016",
  "USGS:04189000:00011:00001",
  "USGS:04189000:00011:00003",
  "USGS:04189000:00011:00007",
  "USGS:04189131:00011:00002",
  "USGS:04189131:00011:00001",
  "USGS:04189174:00011:00002",
  "USGS:04189174:00011:00001",
  "USGS:04189260:00011:00012",
  "USGS:04189260:00011:00002",
  "USGS:04190000:00011:00001",
  "USGS:04190000:00011:00002",
  "USGS:04191500:00011:00009",
  "USGS:04191500:00011:00008",
  "USGS:04192500:00011:00004",
  "USGS:04192500:00011:00003",
  "USGS:04193490:00011:00001",
  "USGS:04193490:00011:00003",
  "USGS:04193490:00011:00004",
  "USGS:04193490:00011:00005",
  "USGS:04193490:00011:00006",
  "USGS:04193500:00011:00001",
  "USGS:04193500:00011:00002",
  "USGS:04195500:00011:00015",
  "USGS:04195500:00011:00001",
  "USGS:04195500:00011:00004",
  "USGS:04195500:00011:00016",
  "USGS:04195500:00011:00017",
  "USGS:04195500:00011:00018",
  "USGS:04195500:00011:00019",
  "USGS:04195820:00011:00004",
  "USGS:04195820:00011:00003",
  "USGS:04196000:00011:00002",
  "USGS:04196000:00011:00001",
  "USGS:04196500:00011:00003",
  "USGS:04196500:00011:00008",
  "USGS:04196800:00011:00002",
  "USGS:04196800:00011:00006",
  "USGS:04197100:00011:00016",
  "USGS:04197100:00011:00009",
  "USGS:04197137:00011:00002",
  "USGS:04197137:00011:00001",
  "USGS:04197170:00011:00001",
  "USGS:04197170:00011:00002",
  "USGS:04198000:00011:00001",
  "USGS:04198000:00011:00020",
  "USGS:04198000:00011:00008",
  "USGS:04199000:00011:00025",
  "USGS:04199000:00011:00024",
  "USGS:04199155:00011:00002",
  "USGS:04199155:00011:00001",
  "USGS:04199500:00011:00001",
  "USGS:04199500:00011:00003",
  "USGS:04199500:00011:00008",
  "USGS:04199500:00011:00004",
  "USGS:04199500:00011:00005",
  "USGS:04199500:00011:00006",
  "USGS:04199500:00011:00020",
  "USGS:04199500:00011:00021",
  "USGS:04200500:00011:00001",
  "USGS:04200500:00011:00002",
  "USGS:04200500:00011:00006",
  "USGS:04200500:00011:00003",
  "USGS:04200500:00011:00019",
  "USGS:04200500:00011:00020",
  "USGS:04200500:00011:00021",
  "USGS:04200500:00011:00022",
  "USGS:04201500:00011:00006",
  "USGS:04201500:00011:00001",
  "USGS:04201500:00011:00004",
  "USGS:04201506:00011:00002",
  "USGS:04201506:00011:00001",
  "USGS:04201515:00011:00007",
  "USGS:04201515:00011:00002",
  "USGS:04201515:00011:00001",
  "USGS:04201526:00011:00011",
  "USGS:04201526:00011:00001",
  "USGS:04202000:00011:00001",
  "USGS:04202000:00011:00007",
  "USGS:04202000:00011:00006",
  "USGS:04206000:00011:00007",
  "USGS:04206000:00011:00006",
  "USGS:04206043:00011:00002",
  "USGS:04206043:00011:00001",
  "USGS:04206212:00011:00002",
  "USGS:04206212:00011:00001",
  "USGS:04206220:00011:00002",
  "USGS:04206220:00011:00001",
  "USGS:04206413:00011:00011",
  "USGS:04206413:00011:00001",
  "USGS:04206416:00011:00002",
  "USGS:04206416:00011:00001",
  "USGS:04206425:00011:00003",
  "USGS:04206425:00011:00002",
  "USGS:04206425:00011:00001",
  "USGS:04206425:00011:00004",
  "USGS:04206448:00011:00002",
  "USGS:04206448:00011:00001",
  "USGS:04207200:00011:00001",
  "USGS:04207200:00011:00004",
  "USGS:04208000:00011:00005",
  "USGS:04208000:00011:00008",
  "USGS:04208000:00011:00007",
  "USGS:04208000:00011:00003",
  "USGS:04208000:00011:00004",
  "USGS:04208000:00011:00006",
  "USGS:04208000:00011:00044",
  "USGS:04208347:00011:00001",
  "USGS:04208460:00011:00002",
  "USGS:04208460:00011:00001",
  "USGS:04208502:00011:00005",
  "USGS:04208504:00011:00001",
  "USGS:04208504:00011:00003",
  "USGS:04208504:00011:00002",
  "USGS:04208700:00011:00011",
  "USGS:04208700:00011:00002",
  "USGS:04208700:00011:00001",
  "USGS:04208700:00011:00012",
  "USGS:04208700:00011:00010",
  "USGS:04208700:00011:00009",
  "USGS:351320080502645:00011:00004",
  "USGS:351331080525945:00011:00004",
  "USGS:351412080541245:00011:00004",
  "USGS:351414080463245:00011:00004",
  "USGS:351455080374445:00011:00004",
  "USGS:351502080512045:00011:00004",
  "USGS:351536080410645:00011:00004",
  "USGS:351540080430045:00011:00001",
  "USGS:351553080562645:00011:00004",
  "USGS:351604080470845:00011:00004",
  "USGS:351609079343701:00011:00001",
  "USGS:351633080493445:00011:00003",
  "USGS:351642080533445:00011:00001",
  "USGS:351709082434101:00011:00001",
  "USGS:351753081011745:00011:00004",
  "USGS:351808082374302:00011:00001",
  "USGS:351812080445545:00011:00001",
  "USGS:351816080564345:00011:00004",
  "USGS:351822081140545:00011:00002",
  "USGS:351849078163901:00011:00001",
  "USGS:351922080540345:00011:00003",
  "USGS:01115190:00011:00004",
  "USGS:01115190:00011:00001",
  "USGS:01115190:00011:00003",
  "USGS:01115265:00011:00003",
  "USGS:01115265:00011:00002",
  "USGS:01115265:00011:00001",
  "USGS:01115265:00011:00004",
  "USGS:01115275:00011:00002",
  "USGS:01115275:00011:00004",
  "USGS:01115275:00011:00001",
  "USGS:01115275:00011:00003",
  "USGS:01115276:00011:00006",
  "USGS:01115276:00011:00002",
  "USGS:01115276:00011:00001",
  "USGS:01115276:00011:00003",
  "USGS:01115280:00011:00002",
  "USGS:01115280:00011:00004",
  "USGS:01115280:00011:00001",
  "USGS:01115280:00011:00003",
  "USGS:01115297:00011:00003",
  "USGS:01115297:00011:00004",
  "USGS:01115297:00011:00001",
  "USGS:01115297:00011:00002",
  "USGS:0208114150:00011:00002",
  "USGS:0208114150:00011:00003",
  "USGS:0208114150:00011:00001",
  "USGS:0208114150:00011:00004",
  "USGS:0208114150:00011:00019",
  "USGS:0208114150:00011:00007",
  "USGS:0208114150:00011:00020",
  "USGS:0208114150:00011:00006",
  "USGS:0208114150:00011:00021",
  "USGS:0208114150:00011:00009",
  "USGS:0208114150:00011:00022",
  "USGS:0208114150:00011:00034",
  "USGS:0208114150:00011:00035",
  "USGS:02081500:00011:00001",
  "USGS:02081500:00011:00002",
  "USGS:02081747:00011:00014",
  "USGS:02081747:00011:00001",
  "USGS:02081747:00011:00002",
  "USGS:02081942:00011:00002",
  "USGS:02081942:00011:00001",
  "USGS:0208250410:00011:00012",
  "USGS:0208250410:00011:00001",
  "USGS:02082585:00011:00014",
  "USGS:02082585:00011:00001",
  "USGS:02082585:00011:00002",
  "USGS:02082770:00011:00001",
  "USGS:02082770:00011:00002",
  "USGS:02082950:00011:00001",
  "USGS:02082950:00011:00002",
  "USGS:02083000:00011:00002",
  "USGS:02083000:00011:00003",
  "USGS:02083500:00011:00002",
  "USGS:02083500:00011:00003",
  "USGS:02084000:00011:00027",
  "USGS:02084000:00011:00021",
  "USGS:02084000:00011:00016",
  "USGS:02084000:00011:00003",
  "USGS:02084160:00011:00002",
  "USGS:02084160:00011:00003",
  "USGS:02084472:00011:00041",
  "USGS:02084557:00011:00002",
  "USGS:02084557:00011:00003",
  "USGS:0208458892:00011:00007",
  "USGS:0208458892:00011:00002",
  "USGS:0208458892:00011:00001",
  "USGS:0208458892:00011:00003",
  "USGS:0208458892:00011:00006",
  "USGS:0208458892:00011:00005",
  "USGS:0208458892:00011:00008",
  "USGS:0208458892:00011:00009",
  "USGS:0208458892:00011:00025",
  "USGS:0208458893:00011:00007",
  "USGS:0208458893:00011:00002",
  "USGS:0208458893:00011:00001",
  "USGS:0208458893:00011:00003",
  "USGS:0208458893:00011:00006",
  "USGS:0208458893:00011:00005",
  "USGS:0208458893:00011:00008",
  "USGS:0208458893:00011:00009",
  "USGS:0208458893:00011:00025",
  "USGS:02085000:00011:00001",
  "USGS:02085000:00011:00002",
  "USGS:02085039:00011:00001",
  "USGS:02085070:00011:00002",
  "USGS:02085070:00011:00003",
  "USGS:0208521324:00011:00002",
  "USGS:0208521324:00011:00001",
  "USGS:0208524090:00011:00002",
  "USGS:0208524090:00011:00001",
  "USGS:0208524975:00011:00002",
  "USGS:0208524975:00011:00001",
  "USGS:02085500:00011:00001",
  "USGS:02085500:00011:00002",
  "USGS:02086500:00011:00002",
  "USGS:02086500:00011:00004",
  "USGS:02086624:00011:00002",
  "USGS:02086624:00011:00004",
  "USGS:0208675010:00011:00002",
  "USGS:0208675010:00011:00001",
  "USGS:02086849:00011:00002",
  "USGS:02086849:00011:00006",
  "USGS:0208700550:00011:00001",
  "USGS:0208706575:00011:00003",
  "USGS:0208706575:00011:00015",
  "USGS:0208706575:00011:00001",
  "USGS:02087182:00011:00001",
  "USGS:02087182:00011:00002",
  "USGS:02087182:00011:00018",
  "USGS:02087182:00011:00004",
  "USGS:02087183:00011:00002",
  "USGS:02087183:00011:00003",
  "USGS:0208726005:00011:00003",
  "USGS:0208726005:00011:00001",
  "USGS:02087275:00011:00003",
  "USGS:02087275:00011:00002",
  "USGS:02087275:00011:00001",
  "USGS:0208731190:00011:00001",
  "USGS:02087322:00011:00014",
  "USGS:02087322:00011:00001",
  "USGS:02087324:00011:00002",
  "USGS:02087324:00011:00001",
  "USGS:0208732534:00011:00003",
  "USGS:0208732534:00011:00002",
  "USGS:0208732534:00011:00001",
  "USGS:0208732885:00011:00002",
  "USGS:0208732885:00011:00003",
  "USGS:0208732885:00011:00005",
  "USGS:0208735012:00011:00016",
  "USGS:0208735012:00011:00005",
  "USGS:0208735012:00011:00001",
  "USGS:02087359:00011:00012",
  "USGS:02087359:00011:00002",
  "USGS:02087359:00011:00001",
  "USGS:02087500:00011:00005",
  "USGS:02087500:00011:00006",
  "USGS:02087570:00011:00003",
  "USGS:02087580:00011:00015",
  "USGS:02087580:00011:00013",
  "USGS:02087580:00011:00001",
  "USGS:02264140:00011:00002",
  "USGS:01116000:00011:00001",
  "USGS:01116000:00011:00003",
  "USGS:01116500:00011:00002",
  "USGS:344544079263701:00011:00001",
  "USGS:345051078012109:00011:00010",
  "USGS:345051078012109:00011:00001",
  "USGS:345609080415102:00011:00001",
  "USGS:345609080415103:00011:00001",
  "USGS:345609080415145:00011:00002",
  "USGS:345809077301408:00011:00001",
  "USGS:345812079313401:00011:00001",
  "USGS:350110080502045:00011:00004",
  "USGS:350314080484945:00011:00001",
  "USGS:350351080454145:00011:00001",
  "USGS:350359080521145:00011:00001",
  "USGS:350623080583801:00011:00001",
  "USGS:350627080410645:00011:00004",
  "USGS:350630080455845:00011:00004",
  "USGS:350635080513245:00011:00004",
  "USGS:350637080475645:00011:00004",
  "USGS:350646080432545:00011:00004",
  "USGS:350657080544945:00011:00003",
  "USGS:350815080460745:00011:00001",
  "USGS:350823080505345:00011:00004",
  "USGS:350842080572801:00011:00001",
  "USGS:350857080383245:00011:00004",
  "USGS:350903081004545:00011:00004",
  "USGS:350947080524945:00011:00002",
  "USGS:351001080495845:00011:00004",
  "USGS:351020079282801:00011:00001",
  "USGS:351023080435745:00011:00001",
  "USGS:351028080385545:00011:00004",
  "USGS:351032080475245:00011:00004",
  "USGS:351104080521845:00011:00004",
  "USGS:351109080412145:00011:00004",
  "USGS:351121083545002:00011:00001",
  "USGS:351124080581245:00011:00002",
  "USGS:351126079301401:00011:00001",
  "USGS:351132079275301:00011:00001",
  "USGS:351132080504145:00011:00001",
  "USGS:351132080562345:00011:00001",
  "USGS:351132080562345:00011:00002",
  "USGS:351134079284901:00011:00001",
  "USGS:351145080371945:00011:00004",
  "USGS:351218079274401:00011:00001",
  "USGS:351218080331345:00011:00004",
  "USGS:351229080460245:00011:00004",
  "USGS:351229080480145:00011:00004",
  "USGS:351247080592745:00011:00004",
  "USGS:351302080412701:00011:00001",
  "USGS:01354330:00011:00001",
  "USGS:01354330:00011:00004",
  "USGS:01354500:00011:00003",
  "USGS:01354500:00011:00004",
  "USGS:01354500:00011:00001",
  "USGS:01355475:00011:00002",
  "USGS:01357500:00011:00003",
  "USGS:01357500:00011:00001",
  "USGS:01357500:00011:00026",
  "USGS:351928080515645:00011:00004",
  "USGS:351943080323145:00011:00002",
  "USGS:351954080493445:00011:00001",
  "USGS:352000080414645:00011:00004",
  "USGS:352003080591245:00011:00003",
  "USGS:352006080462845:00011:00004",
  "USGS:352012081154301:00011:00001",
  "USGS:352012081154302:00011:00001",
  "USGS:352012081154345:00011:00001",
  "USGS:352135080462045:00011:00004",
  "USGS:352155080531145:00011:00003",
  "USGS:352224080500345:00011:00004",
  "USGS:352310080424845:00011:00004",
  "USGS:352315082484401:00011:00001",
  "USGS:352323080551645:00011:00001",
  "USGS:352432080473745:00011:00004",
  "USGS:352440080505045:00011:00004",
  "USGS:352523080535545:00011:00004",
  "USGS:352541080441745:00011:00004",
  "USGS:352555080574445:00011:00004",
  "USGS:352602081014745:00011:00002",
  "USGS:352718080484345:00011:00008",
  "USGS:352750080523545:00011:00003",
  "USGS:352921080473245:00011:00004",
  "USGS:353003080591745:00011:00006",
  "USGS:353014080524945:00011:00004",
  "USGS:353135080524201:00011:00001",
  "USGS:353135080524202:00011:00001",
  "USGS:353135080524203:00011:00001",
  "USGS:01513831:00011:00002",
  "USGS:01513831:00011:00001",
  "USGS:01514000:00011:00002",
  "USGS:01520500:00011:00001",
  "USGS:01520500:00011:00002",
  "USGS:01521000:00011:00002",
  "USGS:01521000:00011:00001",
  "USGS:01521500:00011:00001",
  "USGS:01521500:00011:00015",
  "USGS:01523000:00011:00002",
  "USGS:01523000:00011:00001",
  "USGS:01523500:00011:00001",
  "USGS:01523500:00011:00003",
  "USGS:01524500:00011:00001",
  "USGS:01524500:00011:00005",
  "USGS:01525500:00011:00001",
  "USGS:01525500:00011:00002",
  "USGS:01525981:00011:00002",
  "USGS:01525981:00011:00001",
  "USGS:01526500:00011:00001",
  "USGS:01526500:00011:00002",
  "USGS:01527500:00011:00001",
  "USGS:01527500:00011:00002",
  "USGS:01528320:00011:00001",
  "USGS:01529500:00011:00001",
  "USGS:01529500:00011:00002",
  "USGS:01529950:00011:00001",
  "USGS:01529950:00011:00002",
  "USGS:01530332:00011:00002",
  "USGS:01530332:00011:00001",
  "USGS:02138520:00011:00001",
  "USGS:02140991:00011:00002",
  "USGS:02140991:00011:00001",
  "USGS:02142000:00011:00012",
  "USGS:02142000:00011:00001",
  "USGS:02142000:00011:00002",
  "USGS:02142654:00011:00002",
  "USGS:02142654:00011:00001",
  "USGS:0214265808:00011:00002",
  "USGS:0214265808:00011:00001",
  "USGS:0214266000:00011:00007",
  "USGS:0214266000:00011:00002",
  "USGS:0214266000:00011:00001",
  "USGS:0214266080:00011:00002",
  "USGS:0214266080:00011:00001",
  "USGS:0214269560:00011:00014",
  "USGS:0214269560:00011:00002",
  "USGS:0214269560:00011:00001",
  "USGS:02142900:00011:00001",
  "USGS:02142900:00011:00002",
  "USGS:02142914:00011:00002",
  "USGS:02142914:00011:00001",
  "USGS:0214291555:00011:00002",
  "USGS:0214291555:00011:00001",
  "USGS:0214295600:00011:00002",
  "USGS:0214295600:00011:00001",
  "USGS:0214297160:00011:00002",
  "USGS:0214297160:00011:00001",
  "USGS:02143000:00011:00001",
  "USGS:02143000:00011:00002",
  "USGS:02143040:00011:00017",
  "USGS:02143040:00011:00002",
  "USGS:02143040:00011:00003",
  "USGS:02143500:00011:00002",
  "USGS:02143500:00011:00003",
  "USGS:02144000:00011:00001",
  "USGS:02144000:00011:00002",
  "USGS:02145000:00011:00002",
  "USGS:02145000:00011:00003",
  "USGS:02146211:00011:00002",
  "USGS:02146211:00011:00003",
  "USGS:0214627970:00011:00002",
  "USGS:0214627970:00011:00001",
  "USGS:02146285:00011:00002",
  "USGS:02146285:00011:00001",
  "USGS:02146300:00011:00001",
  "USGS:02146300:00011:00002",
  "USGS:02146315:00011:00002",
  "USGS:02146315:00011:00001",
  "USGS:02146330:00011:00001",
  "USGS:02146348:00011:00002",
  "USGS:02146348:00011:00001",
  "USGS:02146381:00011:00002",
  "USGS:02146381:00011:00001",
  "USGS:0214640410:00011:00001",
  "USGS:02146409:00011:00002",
  "USGS:02146409:00011:00001",
  "USGS:02146420:00011:00001",
  "USGS:0214642825:00011:00002",
  "USGS:0214642825:00011:00001",
  "USGS:0214643770:00011:00001",
  "USGS:0214643820:00011:00002",
  "USGS:0214643820:00011:00001",
  "USGS:0214643860:00011:00001",
  "USGS:02146449:00011:00001",
  "USGS:0214645022:00011:00002",
  "USGS:0214645022:00011:00001",
  "USGS:0214645075:00011:00002",
  "USGS:0214645075:00011:00001",
  "USGS:0214645080:00011:00002",
  "USGS:0214645080:00011:00001",
  "USGS:02146470:00011:00003",
  "USGS:02146470:00011:00004",
  "USGS:02146507:00011:00001",
  "USGS:02146507:00011:00002",
  "USGS:02146530:00011:00002",
  "USGS:02146530:00011:00001",
  "USGS:0214655255:00011:00002",
  "USGS:0214655255:00011:00001",
  "USGS:02146562:00011:00002",
  "USGS:02146562:00011:00001",
  "USGS:0214657975:00011:00002",
  "USGS:0214657975:00011:00001",
  "USGS:02146600:00011:00003",
  "USGS:02146600:00011:00001",
  "USGS:02146600:00011:00002",
  "USGS:02110550:00011:00001",
  "USGS:02146614:00011:00001",
  "USGS:02146670:00011:00001",
  "USGS:0214668150:00011:00001",
  "USGS:02146700:00011:00001",
  "USGS:02146700:00011:00002",
  "USGS:01387420:00011:00001",
  "USGS:01387420:00011:00002",
  "USGS:01387450:00011:00001",
  "USGS:01387450:00011:00002",
  "USGS:01413088:00011:00002",
  "USGS:01413088:00011:00001",
  "USGS:01413398:00011:00002",
  "USGS:01413398:00011:00001",
  "USGS:01413408:00011:00002",
  "USGS:01413408:00011:00003",
  "USGS:01413500:00011:00001",
  "USGS:01413500:00011:00004",
  "USGS:01414000:00011:00001",
  "USGS:01414000:00011:00003",
  "USGS:01414500:00011:00001",
  "USGS:01414500:00011:00003",
  "USGS:01415000:00011:00001",
  "USGS:01415000:00011:00002",
  "USGS:01417000:00011:00001",
  "USGS:01417000:00011:00002",
  "USGS:01417500:00011:00003",
  "USGS:01417500:00011:00007",
  "USGS:01417500:00011:00002",
  "USGS:01420500:00011:00006",
  "USGS:01420500:00011:00002",
  "USGS:02110550:00011:00007",
  "USGS:02110550:00011:00008",
  "USGS:02110550:00011:00009",
  "USGS:02110550:00011:00010",
  "USGS:02110701:00011:00003",
  "USGS:02110701:00011:00013",
  "USGS:02110701:00011:00002",
  "USGS:02110701:00011:00007",
  "USGS:02110701:00011:00020",
  "USGS:02110701:00011:00004",
  "USGS:02110701:00011:00005",
  "USGS:02110701:00011:00010",
  "USGS:02110701:00011:00012",
  "USGS:02110701:00011:00016",
  "USGS:02110704:00011:00013",
  "USGS:02110704:00011:00007",
  "USGS:02110704:00011:00006",
  "USGS:02110704:00011:00014",
  "USGS:02110704:00011:00001",
  "USGS:02110704:00011:00012",
  "USGS:02110704:00011:00027",
  "USGS:02110704:00011:00025",
  "USGS:02110704:00011:00028",
  "USGS:02110725:00011:00001",
  "USGS:02110755:00011:00003",
  "USGS:02110755:00011:00001",
  "USGS:353135080524245:00011:00001",
  "USGS:353219077153801:00011:00002",
  "USGS:354057080362545:00011:00001",
  "USGS:354057080362601:00011:00001",
  "USGS:354133082042201:00011:00001",
  "USGS:354133082042203:00011:00001",
  "USGS:354133082042245:00011:00002",
  "USGS:354302081433201:00011:00001",
  "USGS:354302081433202:00011:00001",
  "USGS:354303080354645:00011:00001",
  "USGS:354353081410545:00011:00002",
  "USGS:354418076463601:00011:00001",
  "USGS:354534082161645:00011:00001",
  "USGS:354616081085101:00011:00001",
  "USGS:354616081085102:00011:00001",
  "USGS:354616081085145:00011:00002",
  "USGS:354822080521501:00011:00001",
  "USGS:354855080134201:00011:00001",
  "USGS:355020078465645:00011:00001",
  "USGS:355031081243202:00011:00001",
  "USGS:355031081243203:00011:00001",
  "USGS:355031081243245:00011:00002",
  "USGS:355037080393045:00011:00009",
  "USGS:355113080230345:00011:00020",
  "USGS:355359080331701:00011:00001",
  "USGS:355511078570745:00011:00001",
  "USGS:355852078572045:00011:00001",
  "USGS:355856078492945:00011:00001",
  "USGS:355944079013401:00011:00001",
  "USGS:360000080444645:00011:00001",
  "USGS:360143078540945:00011:00001",
  "USGS:02100500:00011:00002",
  "USGS:360334078584145:00011:00001",
  "USGS:360419078543145:00011:00001",
  "USGS:360733079552145:00011:00002",
  "USGS:360754080263945:00011:00001",
  "USGS:361011079595401:00011:00001",
  "USGS:361829076163201:00011:00001",
  "USGS:362228075500401:00011:00002",
  "USGS:362228075500401:00011:00003",
  "USGS:362231079410801:00011:00001",
  "USGS:362416080334345:00011:00001",
  "USGS:362954081303800:00011:00001",
  "USGS:363000080584000:00011:00001",
  "USGS:01311875:00011:00019",
  "USGS:01311875:00011:00015",
  "USGS:01311875:00011:00027",
  "USGS:01311875:00011:00016",
  "USGS:01311875:00011:00001",
  "USGS:01311875:00011:00013",
  "USGS:01311875:00011:00018",
  "USGS:01311875:00011:00023",
  "USGS:01311875:00011:00017",
  "USGS:01312000:00011:00001",
  "USGS:01312000:00011:00002",
  "USGS:01314500:00011:00001",
  "USGS:01315000:00011:00001",
  "USGS:01315000:00011:00002",
  "USGS:01315500:00011:00001",
  "USGS:01315500:00011:00002",
  "USGS:01317000:00011:00002",
  "USGS:02088500:00011:00002",
  "USGS:02088500:00011:00003",
  "USGS:02089000:00011:00002",
  "USGS:02089000:00011:00003",
  "USGS:0208925200:00011:00002",
  "USGS:0208925200:00011:00001",
  "USGS:02089500:00011:00002",
  "USGS:02089500:00011:00003",
  "USGS:02090380:00011:00001",
  "USGS:02090380:00011:00002",
  "USGS:02091000:00011:00001",
  "USGS:02091000:00011:00002",
  "USGS:02091500:00011:00002",
  "USGS:02091500:00011:00003",
  "USGS:02091814:00011:00023",
  "USGS:02091814:00011:00018",
  "USGS:0209205053:00011:00001",
  "USGS:02092500:00011:00002",
  "USGS:02092500:00011:00003",
  "USGS:02092554:00011:00003",
  "USGS:02093000:00011:00001",
  "USGS:02093000:00011:00002",
  "USGS:02093800:00011:00012",
  "USGS:02093800:00011:00001",
  "USGS:02093800:00011:00002",
  "USGS:02093877:00011:00002",
  "USGS:02093877:00011:00001",
  "USGS:0209399200:00011:00003",
  "USGS:0209399200:00011:00002",
  "USGS:0209399200:00011:00001",
  "USGS:02094500:00011:00002",
  "USGS:02094500:00011:00003",
  "USGS:02094659:00011:00003",
  "USGS:02094659:00011:00002",
  "USGS:02094659:00011:00001",
  "USGS:02094770:00011:00001",
  "USGS:02094770:00011:00003",
  "USGS:02094770:00011:00002",
  "USGS:02094775:00011:00001",
  "USGS:02094775:00011:00003",
  "USGS:02094775:00011:00002",
  "USGS:02095000:00011:00002",
  "USGS:02095000:00011:00001",
  "USGS:02095000:00011:00003",
  "USGS:02095181:00011:00003",
  "USGS:02095181:00011:00002",
  "USGS:02095181:00011:00001",
  "USGS:02095271:00011:00001",
  "USGS:02095271:00011:00003",
  "USGS:02095271:00011:00002",
  "USGS:02095500:00011:00003",
  "USGS:02095500:00011:00001",
  "USGS:02095500:00011:00002",
  "USGS:0209553650:00011:00001",
  "USGS:0209553650:00011:00003",
  "USGS:0209553650:00011:00002",
  "USGS:02096500:00011:00014",
  "USGS:02096500:00011:00001",
  "USGS:02096500:00011:00002",
  "USGS:02096846:00011:00002",
  "USGS:02096846:00011:00001",
  "USGS:02096960:00011:00002",
  "USGS:02096960:00011:00003",
  "USGS:0209722970:00011:00002",
  "USGS:0209722970:00011:00001",
  "USGS:02097280:00011:00002",
  "USGS:02097280:00011:00001",
  "USGS:02097314:00011:00002",
  "USGS:02097314:00011:00004",
  "USGS:0209734440:00011:00002",
  "USGS:0209734440:00011:00001",
  "USGS:0209741387:00011:00001",
  "USGS:0209741955:00011:00002",
  "USGS:0209741955:00011:00004",
  "USGS:02097464:00011:00002",
  "USGS:02097464:00011:00001",
  "USGS:02097517:00011:00002",
  "USGS:02097517:00011:00004",
  "USGS:0209782609:00011:00011",
  "USGS:0209782609:00011:00001",
  "USGS:02098197:00011:00017",
  "USGS:02098197:00011:00013",
  "USGS:02098197:00011:00010",
  "USGS:02098198:00011:00006",
  "USGS:02098206:00011:00004",
  "USGS:02098206:00011:00007",
  "USGS:02099000:00011:00001",
  "USGS:02099000:00011:00002",
  "USGS:02100500:00011:00003",
  "USGS:0210166029:00011:00002",
  "USGS:0210166029:00011:00001",
  "USGS:02101726:00011:00002",
  "USGS:02101726:00011:00018",
  "USGS:02101726:00011:00001",
  "USGS:02101726:00011:00003",
  "USGS:02101726:00011:00006",
  "USGS:02101726:00011:00005",
  "USGS:02101726:00011:00008",
  "USGS:02101800:00011:00001",
  "USGS:02101800:00011:00002",
  "USGS:02102000:00011:00004",
  "USGS:02102000:00011:00005",
  "USGS:02102192:00011:00001",
  "USGS:02102192:00011:00002",
  "USGS:04273500:00011:00001",
  "USGS:04273500:00011:00002",
  "USGS:04273700:00011:00001",
  "USGS:04273700:00011:00002",
  "USGS:04273800:00011:00002",
  "USGS:04273800:00011:00001",
  "USGS:04275000:00011:00002",
  "USGS:04275500:00011:00001",
  "USGS:04275500:00011:00002",
  "USGS:04276500:00011:00001",
  "USGS:04276500:00011:00002",
  "USGS:04278000:00011:00003",
  "USGS:04279085:00011:00001",
  "USGS:04280450:00011:00002",
  "USGS:0214678175:00011:00001",
  "USGS:0214685800:00011:00002",
  "USGS:0214685800:00011:00001",
  "USGS:02147126:00011:00002",
  "USGS:02147126:00011:00001",
  "USGS:02149000:00011:00001",
  "USGS:02149000:00011:00002",
  "USGS:02150495:00011:00012",
  "USGS:02150495:00011:00002",
  "USGS:02150495:00011:00001",
  "USGS:02151500:00011:00002",
  "USGS:02151500:00011:00003",
  "USGS:02152100:00011:00001",
  "USGS:02152100:00011:00002",
  "USGS:02152474:00011:00002",
  "USGS:02152474:00011:00001",
  "USGS:03161000:00011:00002",
  "USGS:03161000:00011:00003",
  "USGS:03439000:00011:00002",
  "USGS:03439000:00011:00003",
  "USGS:03441000:00011:00001",
  "USGS:03441000:00011:00002",
  "USGS:03443000:00011:00002",
  "USGS:03443000:00011:00003",
  "USGS:03446000:00011:00001",
  "USGS:03446000:00011:00002",
  "USGS:03446000:00011:00003",
  "USGS:03447687:00011:00011",
  "USGS:03447687:00011:00001",
  "USGS:0344894205:00011:00002",
  "USGS:0344894205:00011:00001",
  "USGS:03450000:00011:00002",
  "USGS:03450000:00011:00003",
  "USGS:03451000:00011:00001",
  "USGS:03451000:00011:00002",
  "USGS:03451500:00011:00001",
  "USGS:03451500:00011:00017",
  "USGS:03451500:00011:00002",
  "USGS:03451500:00011:00003",
  "USGS:03453000:00011:00002",
  "USGS:03453000:00011:00003",
  "USGS:03453500:00011:00002",
  "USGS:03453500:00011:00003",
  "USGS:03454500:00011:00002",
  "USGS:03454500:00011:00003",
  "USGS:03455500:00011:00001",
  "USGS:03455500:00011:00002",
  "USGS:03455773:00011:00003",
  "USGS:03455773:00011:00001",
  "USGS:0345577330:00011:00002",
  "USGS:0345577330:00011:00001",
  "USGS:03456100:00011:00001",
  "USGS:03456100:00011:00002",
  "USGS:03456500:00011:00006",
  "USGS:03456500:00011:00002",
  "USGS:03456500:00011:00003",
  "USGS:03456991:00011:00014",
  "USGS:03456991:00011:00002",
  "USGS:03456991:00011:00001",
  "USGS:03459500:00011:00002",
  "USGS:03459500:00011:00003",
  "USGS:03460000:00011:00001",
  "USGS:03460000:00011:00002",
  "USGS:03460000:00011:00003",
  "USGS:03460795:00011:00012",
  "USGS:03460795:00011:00002",
  "USGS:03460795:00011:00001",
  "USGS:03460795:00011:00013",
  "USGS:03460795:00011:00014",
  "USGS:03463300:00011:00002",
  "USGS:03463300:00011:00003",
  "USGS:03479000:00011:00002",
  "USGS:03479000:00011:00003",
  "USGS:03500000:00011:00002",
  "USGS:03500000:00011:00003",
  "USGS:03500240:00011:00001",
  "USGS:03500240:00011:00002",
  "USGS:03501500:00011:00005",
  "USGS:03501500:00011:00001",
  "USGS:03501500:00011:00002",
  "USGS:03501500:00011:00003",
  "USGS:03501500:00011:00006",
  "USGS:03501500:00011:00007",
  "USGS:03501975:00011:00012",
  "USGS:03501975:00011:00002",
  "USGS:03501975:00011:00001",
  "USGS:03501975:00011:00013",
  "USGS:03501975:00011:00014",
  "USGS:03503000:00011:00017",
  "USGS:02129000:00011:00003",
  "USGS:03503000:00011:00001",
  "USGS:03503000:00011:00002",
  "USGS:03504000:00011:00002",
  "USGS:03504000:00011:00003",
  "USGS:03505550:00011:00002",
  "USGS:03505550:00011:00001",
  "USGS:03508050:00011:00002",
  "USGS:03508050:00011:00001",
  "USGS:03510577:00011:00002",
  "USGS:03510577:00011:00001",
  "USGS:03512000:00011:00001",
  "USGS:03512000:00011:00002",
  "USGS:03512000:00011:00025",
  "USGS:03513000:00011:00012",
  "USGS:03513000:00011:00001",
  "USGS:03513000:00011:00002",
  "USGS:0351706800:00011:00012",
  "USGS:0351706800:00011:00002",
  "USGS:0351706800:00011:00001",
  "USGS:03550000:00011:00002",
  "USGS:03550000:00011:00003",
  "USGS:335146078002001:00011:00002",
  "USGS:335146078002001:00011:00003",
  "USGS:335146078002001:00011:00001",
  "USGS:335335078351901:00011:00001",
  "USGS:335629078115406:00011:00001",
  "USGS:335629078115407:00011:00001",
  "USGS:04234000:00011:00001",
  "USGS:04234000:00011:00003",
  "USGS:02111391:00011:00001",
  "USGS:02111391:00011:00012",
  "USGS:0211139110:00011:00002",
  "USGS:0211139110:00011:00001",
  "USGS:02111500:00011:00002",
  "USGS:02111500:00011:00003",
  "USGS:02112000:00011:00002",
  "USGS:02112000:00011:00003",
  "USGS:02112250:00011:00001",
  "USGS:02112250:00011:00002",
  "USGS:02113850:00011:00001",
  "USGS:02113850:00011:00002",
  "USGS:02114450:00011:00001",
  "USGS:02114450:00011:00002",
  "USGS:02115360:00011:00001",
  "USGS:02115360:00011:00002",
  "USGS:02116500:00011:00002",
  "USGS:02116500:00011:00003",
  "USGS:02118000:00011:00002",
  "USGS:02118000:00011:00003",
  "USGS:02118500:00011:00001",
  "USGS:02118500:00011:00002",
  "USGS:02120780:00011:00001",
  "USGS:02120780:00011:00002",
  "USGS:02121500:00011:00004",
  "USGS:02121500:00011:00003",
  "USGS:0212378405:00011:00001",
  "USGS:0212393300:00011:00002",
  "USGS:0212393300:00011:00001",
  "USGS:02124080:00011:00002",
  "USGS:02124080:00011:00001",
  "USGS:0212414900:00011:00002",
  "USGS:0212414900:00011:00001",
  "USGS:0212419274:00011:00002",
  "USGS:0212419274:00011:00001",
  "USGS:02124269:00011:00002",
  "USGS:02124269:00011:00001",
  "USGS:0212427947:00011:00001",
  "USGS:0212430293:00011:00002",
  "USGS:0212430293:00011:00001",
  "USGS:0212430653:00011:00002",
  "USGS:0212430653:00011:00001",
  "USGS:0212433550:00011:00012",
  "USGS:0212433550:00011:00002",
  "USGS:0212433550:00011:00001",
  "USGS:0212466000:00011:00002",
  "USGS:0212466000:00011:00001",
  "USGS:0212467451:00011:00002",
  "USGS:0212467451:00011:00001",
  "USGS:0212467595:00011:00002",
  "USGS:0212467595:00011:00001",
  "USGS:02124692:00011:00002",
  "USGS:02124692:00011:00001",
  "USGS:02126000:00011:00002",
  "USGS:02126000:00011:00003",
  "USGS:02126375:00011:00001",
  "USGS:02128000:00011:00001",
  "USGS:02128000:00011:00002",
  "USGS:02129000:00011:00002",
  "USGS:02132320:00011:00002",
  "USGS:02132320:00011:00001",
  "USGS:02133500:00011:00003",
  "USGS:02133500:00011:00004",
  "USGS:02133624:00011:00002",
  "USGS:02133624:00011:00001",
  "USGS:02134170:00011:00002",
  "USGS:02134170:00011:00001",
  "USGS:02134480:00011:00002",
  "USGS:02134480:00011:00001",
  "USGS:02134500:00011:00002",
  "USGS:02134500:00011:00003",
  "USGS:02234308:00011:00002",
  "USGS:02234308:00011:00001",
  "USGS:421746074180201:00011:00001",
  "USGS:421903074152301:00011:00001",
  "USGS:421932078513701:00011:00001",
  "USGS:421946078274901:00011:00001",
  "USGS:421948074483701:00011:00001",
  "USGS:421948074483702:00011:00001",
  "USGS:422241073274601:00011:00001",
  "USGS:422323076190301:00011:00001",
  "USGS:422445077203301:00011:00001",
  "USGS:422622073410901:00011:00001",
  "USGS:422702079005101:00011:00001",
  "USGS:422710076462901:00011:00001",
  "USGS:422902076475801:00011:00001",
  "USGS:422920076275301:00011:00001",
  "USGS:423143076582601:00011:00001",
  "USGS:01531000:00011:00001",
  "USGS:01531000:00011:00010",
  "USGS:03010820:00011:00012",
  "USGS:03010820:00011:00002",
  "USGS:03010820:00011:00001",
  "USGS:03011020:00011:00030",
  "USGS:03011020:00011:00003",
  "USGS:03011020:00011:00004",
  "USGS:03011020:00011:00018",
  "USGS:03013946:00011:00001",
  "USGS:03014500:00011:00001",
  "USGS:03014500:00011:00016",
  "USGS:04213500:00011:00001",
  "USGS:04213500:00011:00026",
  "USGS:04213500:00011:00009",
  "USGS:04213500:00011:00008",
  "USGS:04213500:00011:00003",
  "USGS:04213500:00011:00022",
  "USGS:04213500:00011:00019",
  "USGS:04213500:00011:00021",
  "USGS:04214500:00011:00006",
  "USGS:04214500:00011:00007",
  "USGS:04215000:00011:00001",
  "USGS:04215000:00011:00006",
  "USGS:04215500:00011:00001",
  "USGS:04215500:00011:00004",
  "USGS:04216418:00011:00001",
  "USGS:04216418:00011:00002",
  "USGS:04217000:00011:00002",
  "USGS:04217000:00011:00006",
  "USGS:04218000:00011:00001",
  "USGS:04218000:00011:00003",
  "USGS:04218518:00011:00001",
  "USGS:04218518:00011:00005",
  "USGS:04220045:00011:00002",
  "USGS:04220045:00011:00001",
  "USGS:0422016550:00011:00002",
  "USGS:0422016550:00011:00001",
  "USGS:04221000:00011:00005",
  "USGS:04221000:00011:00021",
  "USGS:04223000:00011:00005",
  "USGS:04223000:00011:00004",
  "USGS:04224775:00011:00005",
  "USGS:04224775:00011:00017",
  "USGS:04227500:00011:00005",
  "USGS:04227500:00011:00002",
  "USGS:04227500:00011:00025",
  "USGS:04228500:00011:00005",
  "USGS:04228500:00011:00018",
  "USGS:04229500:00011:00004",
  "USGS:04229500:00011:00003",
  "USGS:04230380:00011:00005",
  "USGS:04230380:00011:00016",
  "USGS:04230500:00011:00006",
  "USGS:04230500:00011:00022",
  "USGS:04230500:00011:00034",
  "USGS:04230650:00011:00001",
  "USGS:04231000:00011:00006",
  "USGS:04231000:00011:00017",
  "USGS:04231000:00011:00018",
  "USGS:04231600:00011:00049",
  "USGS:04231600:00011:00003",
  "USGS:04231600:00011:00002",
  "USGS:04231600:00011:00058",
  "USGS:04231600:00011:00050",
  "USGS:04231600:00011:00054",
  "USGS:04231600:00011:00051",
  "USGS:04231600:00011:00053",
  "USGS:04231600:00011:00057",
  "USGS:04232050:00011:00003",
  "USGS:04232050:00011:00002",
  "USGS:04232050:00011:00001",
  "USGS:0423205010:00011:00004",
  "USGS:0423205010:00011:00003",
  "USGS:0423205010:00011:00008",
  "USGS:0423205010:00011:00009",
  "USGS:04232482:00011:00001",
  "USGS:04232482:00011:00003",
  "USGS:04232730:00011:00002",
  "USGS:04232730:00011:00001",
  "USGS:04233255:00011:00002",
  "USGS:04233255:00011:00001",
  "USGS:04233286:00011:00002",
  "USGS:04233286:00011:00001",
  "USGS:04233286:00011:00004",
  "USGS:04233300:00011:00002",
  "USGS:04233300:00011:00001",
  "USGS:04233300:00011:00004",
  "USGS:04233500:00011:00001",
  "USGS:02228500:00011:00001",
  "USGS:02228500:00011:00002",
  "USGS:01318500:00011:00004",
  "USGS:01318500:00011:00002",
  "USGS:01321000:00011:00004",
  "USGS:01321000:00011:00002",
  "USGS:01323500:00011:00002",
  "USGS:01325000:00011:00004",
  "USGS:01325000:00011:00002",
  "USGS:01327500:00011:00002",
  "USGS:01327750:00011:00001",
  "USGS:01327750:00011:00005",
  "USGS:01328770:00011:00001",
  "USGS:01329490:00011:00002",
  "USGS:01329490:00011:00001",
  "USGS:01330000:00011:00006",
  "USGS:01330000:00011:00005",
  "USGS:01330884:00011:00011",
  "USGS:01334500:00011:00001",
  "USGS:01334500:00011:00009",
  "USGS:01335754:00011:00001",
  "USGS:01335754:00011:00004",
  "USGS:01335755:00011:00016",
  "USGS:01335755:00011:00001",
  "USGS:01336000:00011:00002",
  "USGS:01336000:00011:00003",
  "USGS:01338000:00011:00002",
  "USGS:01338000:00011:00001",
  "USGS:01339060:00011:00001",
  "USGS:01339060:00011:00002",
  "USGS:01342602:00011:00001",
  "USGS:01342682:00011:00001",
  "USGS:01342730:00011:00002",
  "USGS:01342743:00011:00001",
  "USGS:01343060:00011:00002",
  "USGS:01343060:00011:00001",
  "USGS:01343403:00011:00002",
  "USGS:01343403:00011:00001",
  "USGS:01343900:00011:00001",
  "USGS:01346000:00011:00001",
  "USGS:01346000:00011:00002",
  "USGS:01347000:00011:00001",
  "USGS:01347000:00011:00002",
  "USGS:01348000:00011:00001",
  "USGS:01348000:00011:00002",
  "USGS:01349000:00011:00002",
  "USGS:01349150:00011:00002",
  "USGS:01349150:00011:00001",
  "USGS:01349527:00011:00001",
  "USGS:01349527:00011:00003",
  "USGS:01349700:00011:00002",
  "USGS:01349700:00011:00003",
  "USGS:01349705:00011:00002",
  "USGS:01349705:00011:00001",
  "USGS:01349711:00011:00002",
  "USGS:01349711:00011:00001",
  "USGS:01349810:00011:00002",
  "USGS:01349810:00011:00001",
  "USGS:01349950:00011:00002",
  "USGS:01349950:00011:00001",
  "USGS:01350000:00011:00001",
  "USGS:01350000:00011:00002",
  "USGS:01350000:00011:00014",
  "USGS:01350035:00011:00002",
  "USGS:01350035:00011:00001",
  "USGS:01350080:00011:00002",
  "USGS:01350080:00011:00001",
  "USGS:01350080:00011:00012",
  "USGS:01350100:00011:00001",
  "USGS:01350100:00011:00013",
  "USGS:01350101:00011:00001",
  "USGS:01350101:00011:00002",
  "USGS:01350101:00011:00003",
  "USGS:01350120:00011:00001",
  "USGS:01350120:00011:00002",
  "USGS:01350120:00011:00012",
  "USGS:01350140:00011:00001",
  "USGS:01350140:00011:00003",
  "USGS:01350180:00011:00002",
  "USGS:01350180:00011:00004",
  "USGS:01350355:00011:00002",
  "USGS:01350355:00011:00001",
  "USGS:01350355:00011:00003",
  "USGS:01351500:00011:00002",
  "USGS:01351500:00011:00003",
  "USGS:01351500:00011:00015",
  "USGS:02236125:00011:00007",
  "USGS:02236125:00011:00006",
  "USGS:02236125:00011:00001",
  "USGS:02236125:00011:00008",
  "USGS:02236125:00011:00009",
  "USGS:02236125:00011:00014",
  "USGS:02236125:00011:00010",
  "USGS:02236125:00011:00012",
  "USGS:0423401815:00011:00002",
  "USGS:0423401815:00011:00001",
  "USGS:0423406130:00011:00001",
  "USGS:04234254:00011:00001",
  "USGS:04235000:00011:00001",
  "USGS:04235000:00011:00003",
  "USGS:04235250:00011:00001",
  "USGS:04235250:00011:00003",
  "USGS:04235299:00011:00001",
  "USGS:04235299:00011:00002",
  "USGS:04235396:00011:00002",
  "USGS:04235440:00011:00002",
  "USGS:04235440:00011:00001",
  "USGS:04235600:00011:00022",
  "USGS:04235600:00011:00021",
  "USGS:04236800:00011:00002",
  "USGS:04237500:00011:00006",
  "USGS:04237500:00011:00011",
  "USGS:04237962:00011:00024",
  "USGS:04237962:00011:00002",
  "USGS:04237962:00011:00001",
  "USGS:04239000:00011:00001",
  "USGS:04239000:00011:00003",
  "USGS:04240010:00011:00001",
  "USGS:04240010:00011:00002",
  "USGS:04240100:00011:00001",
  "USGS:04240100:00011:00002",
  "USGS:04240105:00011:00020",
  "USGS:04240105:00011:00022",
  "USGS:04240120:00011:00021",
  "USGS:04240120:00011:00023",
  "USGS:04240300:00011:00001",
  "USGS:04240300:00011:00002",
  "USGS:04240495:00011:00001",
  "USGS:04242500:00011:00002",
  "USGS:04242500:00011:00005",
  "USGS:04242640:00011:00002",
  "USGS:04243500:00011:00001",
  "USGS:04243500:00011:00003",
  "USGS:04243783:00011:00002",
  "USGS:04244000:00011:00002",
  "USGS:04245840:00011:00002",
  "USGS:04245840:00011:00004",
  "USGS:04247000:00011:00024",
  "USGS:04247000:00011:00008",
  "USGS:04247055:00011:00002",
  "USGS:04247055:00011:00001",
  "USGS:04249000:00011:00001",
  "USGS:04249000:00011:00002",
  "USGS:04249000:00011:00007",
  "USGS:04249000:00011:00003",
  "USGS:04249000:00011:00028",
  "USGS:04249000:00011:00025",
  "USGS:04249000:00011:00027",
  "USGS:04249200:00011:00002",
  "USGS:04249200:00011:00001",
  "USGS:04250200:00011:00002",
  "USGS:04250200:00011:00001",
  "USGS:04250750:00011:00002",
  "USGS:04250750:00011:00003",
  "USGS:04252500:00011:00004",
  "USGS:04252500:00011:00002",
  "USGS:04253300:00011:00002",
  "USGS:04254500:00011:00002",
  "USGS:04256000:00011:00002",
  "USGS:04256000:00011:00004",
  "USGS:04256500:00011:00002",
  "USGS:04258000:00011:00001",
  "USGS:04258000:00011:00002",
  "USGS:04260500:00011:00005",
  "USGS:04260500:00011:00002",
  "USGS:04262000:00011:00001",
  "USGS:04262000:00011:00002",
  "USGS:04262500:00011:00001",
  "USGS:04262500:00011:00003",
  "USGS:04263000:00011:00002",
  "USGS:04263000:00011:00003",
  "USGS:04265432:00011:00002",
  "USGS:04265432:00011:00001",
  "USGS:04266500:00011:00001",
  "USGS:04266500:00011:00003",
  "USGS:04267500:00011:00001",
  "USGS:04267500:00011:00002",
  "USGS:04268000:00011:00002",
  "USGS:04268000:00011:00003",
  "USGS:04268800:00011:00001",
  "USGS:04268800:00011:00003",
  "USGS:04269000:00011:00002",
  "USGS:04269000:00011:00003",
  "USGS:04270200:00011:00001",
  "USGS:04270200:00011:00002",
  "USGS:04271500:00011:00001",
  "USGS:04271500:00011:00003",
  "USGS:02270500:00011:00001",
  "USGS:02270500:00011:00002",
  "USGS:02271500:00011:00001",
  "USGS:02271500:00011:00002",
  "USGS:02272650:00011:00002",
  "USGS:02272650:00011:00001",
  "USGS:02272676:00011:00002",
  "USGS:02272676:00011:00001",
  "USGS:02273230:00011:00002",
  "USGS:02273230:00011:00001",
  "USGS:02273630:00011:00002",
  "USGS:02273630:00011:00001",
  "USGS:02274005:00011:00002",
  "USGS:02274005:00011:00001",
  "USGS:02274010:00011:00002",
  "USGS:02274010:00011:00001",
  "USGS:02274325:00011:00002",
  "USGS:02274325:00011:00001",
  "USGS:02274490:00011:00002",
  "USGS:02274490:00011:00001",
  "USGS:02274505:00011:00002",
  "USGS:02274505:00011:00001",
  "USGS:02275197:00011:00002",
  "USGS:02275197:00011:00001",
  "USGS:02276877:00011:00050",
  "USGS:02276877:00011:00047",
  "USGS:02276877:00011:00003",
  "USGS:02277100:00011:00005",
  "USGS:02277100:00011:00007",
  "USGS:01421000:00011:00003",
  "USGS:01421000:00011:00002",
  "USGS:01421000:00011:00007",
  "USGS:01421610:00011:00002",
  "USGS:01421610:00011:00001",
  "USGS:01421618:00011:00002",
  "USGS:01421618:00011:00001",
  "USGS:01421900:00011:00002",
  "USGS:01421900:00011:00003",
  "USGS:01422500:00011:00001",
  "USGS:01422500:00011:00002",
  "USGS:01423000:00011:00001",
  "USGS:01423000:00011:00002",
  "USGS:0142400103:00011:00002",
  "USGS:0142400103:00011:00001",
  "USGS:01425000:00011:00004",
  "USGS:01425000:00011:00002",
  "USGS:01425000:00011:00003",
  "USGS:01426500:00011:00003",
  "USGS:01426500:00011:00007",
  "USGS:01426500:00011:00002",
  "USGS:01427000:00011:00001",
  "USGS:01427500:00011:00004",
  "USGS:01428500:00011:00001",
  "USGS:01428500:00011:00002",
  "USGS:01428500:00011:00006",
  "USGS:01432900:00011:00002",
  "USGS:01432900:00011:00001",
  "USGS:01433500:00011:00003",
  "USGS:01433500:00011:00001",
  "USGS:01433500:00011:00002",
  "USGS:01433500:00011:00004",
  "USGS:01433500:00011:00006",
  "USGS:01433500:00011:00007",
  "USGS:01433500:00011:00005",
  "USGS:01434017:00011:00002",
  "USGS:01434017:00011:00001",
  "USGS:01434025:00011:00001",
  "USGS:01434025:00011:00006",
  "USGS:01434498:00011:00002",
  "USGS:01434498:00011:00012",
  "USGS:01435000:00011:00016",
  "USGS:01435000:00011:00001",
  "USGS:01435000:00011:00017",
  "USGS:01436000:00011:00001",
  "USGS:01436000:00011:00002",
  "USGS:01436690:00011:00005",
  "USGS:01436690:00011:00002",
  "USGS:01436690:00011:00003",
  "USGS:01437500:00011:00002",
  "USGS:01437500:00011:00003",
  "USGS:01499500:00011:00002",
  "USGS:01499500:00011:00001",
  "USGS:01500000:00011:00001",
  "USGS:01500000:00011:00002",
  "USGS:01500500:00011:00002",
  "USGS:01502500:00011:00001",
  "USGS:01502500:00011:00002",
  "USGS:01502632:00011:00002",
  "USGS:01502632:00011:00001",
  "USGS:01502731:00011:00002",
  "USGS:01502731:00011:00001",
  "USGS:01503000:00011:00003",
  "USGS:01503000:00011:00001",
  "USGS:01503000:00011:00002",
  "USGS:01503000:00011:00017",
  "USGS:01503500:00011:00001",
  "USGS:01505000:00011:00001",
  "USGS:01505000:00011:00002",
  "USGS:01505810:00011:00002",
  "USGS:01505810:00011:00001",
  "USGS:01507000:00011:00004",
  "USGS:01507000:00011:00001",
  "USGS:01507000:00011:00002",
  "USGS:01507000:00011:00019",
  "USGS:01509000:00011:00015",
  "USGS:01509000:00011:00001",
  "USGS:01509000:00011:00002",
  "USGS:01509520:00011:00001",
  "USGS:01510000:00011:00003",
  "USGS:01510000:00011:00001",
  "USGS:01510000:00011:00002",
  "USGS:01511500:00011:00002",
  "USGS:01512500:00011:00001",
  "USGS:01512500:00011:00002",
  "USGS:01513500:00011:00001",
  "USGS:01513500:00011:00002",
  "USGS:02249500:00011:00001",
  "USGS:02249500:00011:00002",
  "USGS:02249500:00011:00004",
  "USGS:02249500:00011:00005",
  "USGS:04280450:00011:00003",
  "USGS:04295000:00011:00003",
  "USGS:403547074090801:00011:00001",
  "USGS:403827074060101:00011:00001",
  "USGS:404205073474101:00011:00001",
  "USGS:404505073131501:00011:00001",
  "USGS:404553073351201:00011:00001",
  "USGS:405149072532201:00011:00001",
  "USGS:405249073010701:00011:00001",
  "USGS:405743072425701:00011:00001",
  "USGS:405756072173502:00011:00001",
  "USGS:405830072331502:00011:00001",
  "USGS:405925072165601:00011:00001",
  "USGS:410254072275201:00011:00005",
  "USGS:410254072275201:00011:00002",
  "USGS:410254072275201:00011:00003",
  "USGS:410254072275201:00011:00001",
  "USGS:410254072275201:00011:00004",
  "USGS:410518074020300:00011:00001",
  "USGS:410828074065801:00011:00001",
  "USGS:410853073554001:00011:00001",
  "USGS:411405074141501:00011:00002",
  "USGS:411421073481202:00011:00001",
  "USGS:411802073593001:00011:00001",
  "USGS:412149073445601:00011:00001",
  "USGS:412637074362301:00011:00001",
  "USGS:412714073331301:00011:00001",
  "USGS:413428074085701:00011:00001",
  "USGS:423530074191701:00011:00001",
  "USGS:414128073475201:00011:00001",
  "USGS:414429074052001:00011:00001",
  "USGS:414525074360601:00011:00001",
  "USGS:414737073563301:00011:00001",
  "USGS:414948074035001:00011:00001",
  "USGS:420326079295801:00011:00001",
  "USGS:420530078445201:00011:00001",
  "USGS:420703079442501:00011:00001",
  "USGS:420828076484601:00011:00001",
  "USGS:421138075511301:00011:00001",
  "USGS:421157075535401:00011:00001",
  "USGS:421213076313301:00011:00001",
  "USGS:421429079295601:00011:00001",
  "USGS:421511079161701:00011:00001",
  "USGS:421512077472801:00011:00001",
  "USGS:421544078021301:00011:00001",
  "USGS:421556075281602:00011:00001",
  "USGS:421734079063801:00011:00001",
  "USGS:02299230:00011:00005",
  "USGS:02299230:00011:00006",
  "USGS:02299230:00011:00001",
  "USGS:02299230:00011:00003",
  "USGS:02299230:00011:00004",
  "USGS:02299410:00011:00001",
  "USGS:02299410:00011:00002",
  "USGS:02299450:00011:00003",
  "USGS:02299450:00011:00002",
  "USGS:02299450:00011:00001",
  "USGS:423534073423401:00011:00001",
  "USGS:423743078070802:00011:00002",
  "USGS:423827076035901:00011:00001",
  "USGS:424017074301501:00011:00001",
  "USGS:424115073495301:00011:00001",
  "USGS:424136075025101:00011:00001",
  "USGS:424158076251901:00011:00001",
  "USGS:424311073423901:00011:00001",
  "USGS:424347076530201:00011:00001",
  "USGS:424347076530202:00011:00001",
  "USGS:424452076081902:00011:00001",
  "USGS:424859073585501:00011:00001",
  "USGS:425048073472501:00011:00001",
  "USGS:425448076350002:00011:00001",
  "USGS:425511074254001:00011:00001",
  "USGS:425704078360601:00011:00001",
  "USGS:425803077151201:00011:00001",
  "USGS:425821076461301:00011:00001",
  "USGS:425833077503901:00011:00001",
  "USGS:425840077133901:00011:00001",
  "USGS:425846075504501:00011:00001",
  "USGS:425913078085501:00011:00001",
  "USGS:430056075354102:00011:00001",
  "USGS:430121074523001:00011:00001",
  "USGS:430146078101301:00011:00001",
  "USGS:430243076180401:00011:00001",
  "USGS:430243076180402:00011:00001",
  "USGS:430252077283402:00011:00001",
  "USGS:430311077051501:00011:00001",
  "USGS:430327073475401:00011:00001",
  "USGS:430739078502701:00011:00001",
  "USGS:430924078241301:00011:00001",
  "USGS:431030073192101:00011:00001",
  "USGS:02291669:00011:00002",
  "USGS:02291669:00011:00001",
  "USGS:02291673:00011:00002",
  "USGS:02291673:00011:00001",
  "USGS:02291710:00011:00001",
  "USGS:02291710:00011:00030",
  "USGS:02292010:00011:00004",
  "USGS:02292010:00011:00012",
  "USGS:02292010:00011:00013",
  "USGS:02292010:00011:00006",
  "USGS:02292010:00011:00001",
  "USGS:02292900:00011:00049",
  "USGS:02292900:00011:00003",
  "USGS:02292900:00011:00041",
  "USGS:02292900:00011:00047",
  "USGS:02292900:00011:00048",
  "USGS:02292900:00011:00051",
  "USGS:02292900:00011:00050",
  "USGS:02293230:00011:00002",
  "USGS:02293230:00011:00001",
  "USGS:02293254:00011:00009",
  "USGS:02293254:00011:00005",
  "USGS:02293254:00011:00001",
  "USGS:01116500:00011:00005",
  "USGS:01116905:00011:00001",
  "USGS:01116905:00011:00002",
  "USGS:01117000:00011:00002",
  "USGS:01117000:00011:00004",
  "USGS:01117350:00011:00002",
  "USGS:01117350:00011:00005",
  "USGS:01117370:00011:00002",
  "USGS:01117370:00011:00001",
  "USGS:01117420:00011:00002",
  "USGS:01117420:00011:00005",
  "USGS:01117430:00011:00002",
  "USGS:01117430:00011:00001",
  "USGS:01117468:00011:00002",
  "USGS:01117468:00011:00005",
  "USGS:01117500:00011:00001",
  "USGS:01117500:00011:00004",
  "USGS:01117800:00011:00001",
  "USGS:01117800:00011:00002",
  "USGS:01118000:00011:00002",
  "USGS:01118000:00011:00004",
  "USGS:01118500:00011:00002",
  "USGS:01118500:00011:00003",
  "USGS:01200000:00011:00014",
  "USGS:01200000:00011:00016",
  "USGS:01200000:00011:00002",
  "USGS:01200000:00011:00003",
  "USGS:01302020:00011:00002",
  "USGS:01302020:00011:00001",
  "USGS:01302250:00011:00008",
  "USGS:01302250:00011:00005",
  "USGS:01302250:00011:00006",
  "USGS:01302250:00011:00001",
  "USGS:01302250:00011:00004",
  "USGS:01302250:00011:00007",
  "USGS:01302600:00011:00001",
  "USGS:01302600:00011:00004",
  "USGS:01302845:00011:00008",
  "USGS:01302845:00011:00005",
  "USGS:01302845:00011:00006",
  "USGS:01302845:00011:00001",
  "USGS:01302845:00011:00004",
  "USGS:01302845:00011:00007",
  "USGS:01303500:00011:00001",
  "USGS:01303500:00011:00002",
  "USGS:01304000:00011:00002",
  "USGS:01304000:00011:00004",
  "USGS:01304057:00011:00026",
  "USGS:01304057:00011:00018",
  "USGS:01304057:00011:00019",
  "USGS:01304057:00011:00022",
  "USGS:01304057:00011:00024",
  "USGS:01304057:00011:00001",
  "USGS:01304057:00011:00004",
  "USGS:01304057:00011:00025",
  "USGS:01304057:00011:00021",
  "USGS:01304200:00011:00027",
  "USGS:01304200:00011:00019",
  "USGS:01304200:00011:00020",
  "USGS:01304200:00011:00023",
  "USGS:01304200:00011:00025",
  "USGS:01304200:00011:00001",
  "USGS:01304200:00011:00005",
  "USGS:01304200:00011:00026",
  "USGS:01304200:00011:00022",
  "USGS:01304200:00011:00030",
  "USGS:01304250:00011:00001",
  "USGS:01304500:00011:00002",
  "USGS:01304500:00011:00004",
  "USGS:01304562:00011:00027",
  "USGS:01304562:00011:00019",
  "USGS:01304562:00011:00020",
  "USGS:01304562:00011:00023",
  "USGS:01304562:00011:00026",
  "USGS:01304562:00011:00001",
  "USGS:01304562:00011:00005",
  "USGS:01304562:00011:00025",
  "USGS:01304562:00011:00022",
  "USGS:01304562:00011:00030",
  "USGS:01304705:00011:00001",
  "USGS:01306460:00011:00001",
  "USGS:01306460:00011:00002",
  "USGS:01308500:00011:00001",
  "USGS:01308500:00011:00002",
  "USGS:01309225:00011:00001",
  "USGS:01309225:00011:00013",
  "USGS:01309500:00011:00003",
  "USGS:01309500:00011:00004",
  "USGS:01309950:00011:00001",
  "USGS:01309950:00011:00002",
  "USGS:01310521:00011:00001",
  "USGS:01310521:00011:00011",
  "USGS:01310740:00011:00035",
  "USGS:01310740:00011:00006",
  "USGS:01310740:00011:00005",
  "USGS:01310740:00011:00004",
  "USGS:01310740:00011:00002",
  "USGS:01310740:00011:00007",
  "USGS:01310740:00011:00028",
  "USGS:01310740:00011:00031",
  "USGS:01310740:00011:00010",
  "USGS:01310740:00011:00011",
  "USGS:01310740:00011:00036",
  "USGS:01310740:00011:00027",
  "USGS:01310740:00011:00001",
  "USGS:01310740:00011:00012",
  "USGS:01310740:00011:00034",
  "USGS:01310740:00011:00008",
  "USGS:01310740:00011:00003",
  "USGS:01310740:00011:00030",
  "USGS:01311143:00011:00027",
  "USGS:01311143:00011:00019",
  "USGS:01311143:00011:00020",
  "USGS:01311143:00011:00023",
  "USGS:01311143:00011:00033",
  "USGS:01311143:00011:00035",
  "USGS:01311143:00011:00026",
  "USGS:01311143:00011:00001",
  "USGS:01311143:00011:00005",
  "USGS:01311143:00011:00025",
  "USGS:01311143:00011:00034",
  "USGS:01311143:00011:00022",
  "USGS:01311143:00011:00030",
  "USGS:01311145:00011:00001",
  "USGS:01311145:00011:00013",
  "USGS:01311500:00011:00001",
  "USGS:01311500:00011:00002",
  "USGS:01311850:00011:00001",
  "USGS:01311850:00011:00013",
  "USGS:05049995:00011:00001",
  "USGS:05049995:00011:00002",
  "USGS:05050000:00011:00015",
  "USGS:05050000:00011:00014",
  "USGS:05290000:00011:00001",
  "USGS:05290000:00011:00002",
  "USGS:05291000:00011:00008",
  "USGS:05291000:00011:00007",
  "USGS:06334500:00011:00010",
  "USGS:06334500:00011:00002",
  "USGS:06334500:00011:00008",
  "USGS:06354882:00011:00015",
  "USGS:06354882:00011:00001",
  "USGS:06354882:00011:00003",
  "USGS:06355500:00011:00006",
  "USGS:06355500:00011:00001",
  "USGS:06355500:00011:00004",
  "USGS:412154071462901:00011:00001",
  "USGS:412844071422802:00011:00001",
  "USGS:412918071321001:00011:00001",
  "USGS:412932071374302:00011:00001",
  "USGS:413252071323601:00011:00001",
  "USGS:413358071433801:00011:00001",
  "USGS:01358000:00011:00028",
  "USGS:01358000:00011:00002",
  "USGS:01359139:00011:00005",
  "USGS:01359139:00011:00006",
  "USGS:01360640:00011:00002",
  "USGS:01360640:00011:00003",
  "USGS:01361000:00011:00001",
  "USGS:01361000:00011:00002",
  "USGS:01362090:00011:00003",
  "USGS:01362090:00011:00001",
  "USGS:01362090:00011:00004",
  "USGS:01362090:00011:00015",
  "USGS:013621955:00011:00002",
  "USGS:013621955:00011:00001",
  "USGS:01362200:00011:00002",
  "USGS:01362200:00011:00004",
  "USGS:01362230:00011:00005",
  "USGS:01362230:00011:00002",
  "USGS:01362230:00011:00003",
  "USGS:0136230002:00011:00002",
  "USGS:0136230002:00011:00001",
  "USGS:01362332:00011:00003",
  "USGS:01362342:00011:00002",
  "USGS:01362342:00011:00001",
  "USGS:01362350:00011:00003",
  "USGS:01362356:00011:00003",
  "USGS:01362357:00011:00004",
  "USGS:01362370:00011:00002",
  "USGS:01362370:00011:00001",
  "USGS:01362370:00011:00015",
  "USGS:01362497:00011:00002",
  "USGS:01362497:00011:00001",
  "USGS:01362500:00011:00005",
  "USGS:01362500:00011:00001",
  "USGS:01362500:00011:00006",
  "USGS:01363382:00011:00002",
  "USGS:01363382:00011:00001",
  "USGS:01363556:00011:00002",
  "USGS:01363556:00011:00001",
  "USGS:01363556:00011:00003",
  "USGS:01364500:00011:00001",
  "USGS:01364500:00011:00002",
  "USGS:01364500:00011:00020",
  "USGS:01365000:00011:00001",
  "USGS:01365000:00011:00003",
  "USGS:01365500:00011:00004",
  "USGS:01365500:00011:00003",
  "USGS:01367500:00011:00001",
  "USGS:01367500:00011:00005",
  "USGS:01371500:00011:00002",
  "USGS:01371500:00011:00003",
  "USGS:01372007:00011:00003",
  "USGS:01372007:00011:00004",
  "USGS:01372007:00011:00001",
  "USGS:01372007:00011:00005",
  "USGS:01372043:00011:00003",
  "USGS:01372043:00011:00004",
  "USGS:01372058:00011:00001",
  "USGS:01372058:00011:00048",
  "USGS:01372058:00011:00037",
  "USGS:01372058:00011:00080",
  "USGS:01372058:00011:00007",
  "USGS:01372058:00011:00002",
  "USGS:01372058:00011:00072",
  "USGS:01372500:00011:00002",
  "USGS:01372500:00011:00003",
  "USGS:0137449480:00011:00002",
  "USGS:0137449480:00011:00003",
  "USGS:01374505:00011:00002",
  "USGS:01374505:00011:00003",
  "USGS:01374531:00011:00005",
  "USGS:01374531:00011:00019",
  "USGS:01374559:00011:00002",
  "USGS:01374559:00011:00003",
  "USGS:01374581:00011:00002",
  "USGS:01374581:00011:00001",
  "USGS:01374598:00011:00002",
  "USGS:01374598:00011:00001",
  "USGS:0137462010:00011:00002",
  "USGS:0137462010:00011:00003",
  "USGS:01374701:00011:00002",
  "USGS:01374701:00011:00003",
  "USGS:01374781:00011:00002",
  "USGS:01374781:00011:00001",
  "USGS:01374821:00011:00002",
  "USGS:01374821:00011:00003",
  "USGS:01374890:00011:00002",
  "USGS:01374890:00011:00003",
  "USGS:01374901:00011:00002",
  "USGS:01374901:00011:00003",
  "USGS:01374930:00011:00002",
  "USGS:01374930:00011:00003",
  "USGS:01374941:00011:00002",
  "USGS:01374941:00011:00003",
  "USGS:01375000:00011:00001",
  "USGS:01375000:00011:00002",
  "USGS:01376269:00011:00001",
  "USGS:01376269:00011:00003",
  "USGS:01376269:00011:00002",
  "USGS:01376800:00011:00001",
  "USGS:01376800:00011:00002",
  "USGS:01387400:00011:00001",
  "USGS:01387400:00011:00002",
  "USGS:02310288:00011:00001",
  "USGS:02310300:00011:00001",
  "USGS:02310300:00011:00002",
  "USGS:02310300:00011:00016",
  "USGS:02310308:00011:00003",
  "USGS:02310308:00011:00001",
  "USGS:02310308:00011:00002",
  "USGS:02310368:00011:00011",
  "USGS:02310368:00011:00001",
  "USGS:02310525:00011:00017",
  "USGS:02310650:00011:00026",
  "USGS:02310650:00011:00022",
  "USGS:02310650:00011:00021",
  "USGS:02310650:00011:00027",
  "USGS:02310650:00011:00029",
  "USGS:02310663:00011:00011",
  "USGS:02310663:00011:00013",
  "USGS:02277100:00011:00001",
  "USGS:02277100:00011:00026",
  "USGS:02277100:00011:00027",
  "USGS:02277100:00011:00028",
  "USGS:02277100:00011:00029",
  "USGS:02277110:00011:00005",
  "USGS:02277110:00011:00007",
  "USGS:02277110:00011:00001",
  "USGS:02277110:00011:00028",
  "USGS:02277110:00011:00029",
  "USGS:02277110:00011:00030",
  "USGS:02277110:00011:00031",
  "USGS:02277110:00011:00008",
  "USGS:02277600:00011:00001",
  "USGS:02277600:00011:00002",
  "USGS:02277600:00011:00004",
  "USGS:02277602:00011:00001",
  "USGS:02277602:00011:00002",
  "USGS:02280500:00011:00035",
  "USGS:02280500:00011:00021",
  "USGS:02280500:00011:00022",
  "USGS:02281200:00011:00046",
  "USGS:02281200:00011:00001",
  "USGS:02281200:00011:00002",
  "USGS:02281200:00011:00007",
  "USGS:02283500:00011:00022",
  "USGS:02283500:00011:00023",
  "USGS:02286400:00011:00041",
  "USGS:02286400:00011:00002",
  "USGS:02286400:00011:00003",
  "USGS:02287497:00011:00026",
  "USGS:02287497:00011:00029",
  "USGS:02287497:00011:00030",
  "USGS:02288800:00011:00003",
  "USGS:02288800:00011:00004",
  "USGS:02288800:00011:00015",
  "USGS:02288900:00011:00001",
  "USGS:02288900:00011:00003",
  "USGS:02289019:00011:00016",
  "USGS:02289019:00011:00024",
  "USGS:02289019:00011:00007",
  "USGS:02289019:00011:00008",
  "USGS:02289035:00011:00003",
  "USGS:02289035:00011:00002",
  "USGS:02289035:00011:00028",
  "USGS:02289035:00011:00027",
  "USGS:02289041:00011:00003",
  "USGS:02289041:00011:00015",
  "USGS:02289041:00011:00024",
  "USGS:02289041:00011:00025",
  "USGS:02289060:00011:00002",
  "USGS:02289060:00011:00012",
  "USGS:02289500:00011:00003",
  "USGS:02289500:00011:00001",
  "USGS:02289500:00011:00002",
  "USGS:02289500:00011:00008",
  "USGS:022907085:00011:00003",
  "USGS:022907085:00011:00001",
  "USGS:022907085:00011:00002",
  "USGS:022907085:00011:00004",
  "USGS:022907647:00011:00026",
  "USGS:022907647:00011:00031",
  "USGS:022907647:00011:00001",
  "USGS:02290765:00011:00025",
  "USGS:02290765:00011:00030",
  "USGS:02290765:00011:00001",
  "USGS:02290766:00011:00020",
  "USGS:02290766:00011:00015",
  "USGS:02290766:00011:00001",
  "USGS:02290767:00011:00048",
  "USGS:02290767:00011:00016",
  "USGS:02290767:00011:00001",
  "USGS:02290768:00011:00021",
  "USGS:02290768:00011:00015",
  "USGS:02290768:00011:00001",
  "USGS:02290769:00011:00034",
  "USGS:02290769:00011:00001",
  "USGS:02290769:00011:00007",
  "USGS:02290769:00011:00012",
  "USGS:022908205:00011:00009",
  "USGS:022908205:00011:00051",
  "USGS:022908205:00011:00060",
  "USGS:022908205:00011:00001",
  "USGS:022908205:00011:00053",
  "USGS:022908205:00011:00026",
  "USGS:022908205:00011:00007",
  "USGS:022908205:00011:00056",
  "USGS:022908295:00011:00007",
  "USGS:022908295:00011:00027",
  "USGS:022908295:00011:00041",
  "USGS:022908295:00011:00023",
  "USGS:022908295:00011:00039",
  "USGS:022908295:00011:00009",
  "USGS:022908295:00011:00010",
  "USGS:02290878:00011:00008",
  "USGS:02290878:00011:00004",
  "USGS:02290878:00011:00001",
  "USGS:02290878:00011:00006",
  "USGS:02290878:00011:00023",
  "USGS:02290888:00011:00008",
  "USGS:02290888:00011:00004",
  "USGS:02290888:00011:00001",
  "USGS:02290888:00011:00006",
  "USGS:02290888:00011:00026",
  "USGS:02290918:00011:00009",
  "USGS:02290918:00011:00002",
  "USGS:02290918:00011:00004",
  "USGS:02290918:00011:00021",
  "USGS:02290918:00011:00007",
  "USGS:02290918:00011:00027",
  "USGS:02290928:00011:00003",
  "USGS:02290928:00011:00001",
  "USGS:02290928:00011:00004",
  "USGS:02290928:00011:00002",
  "USGS:02290930:00011:00003",
  "USGS:02290930:00011:00001",
  "USGS:02290930:00011:00002",
  "USGS:02290942:00011:00003",
  "USGS:02290942:00011:00015",
  "USGS:02290942:00011:00004",
  "USGS:02290942:00011:00001",
  "USGS:02290942:00011:00002",
  "USGS:02290942:00011:00005",
  "USGS:02291001:00011:00001",
  "USGS:02291001:00011:00002",
  "USGS:02291200:00011:00002",
  "USGS:02291500:00011:00001",
  "USGS:02291500:00011:00002",
  "USGS:02291524:00011:00002",
  "USGS:02291524:00011:00001",
  "USGS:02291580:00011:00002",
  "USGS:02291580:00011:00001",
  "USGS:02291597:00011:00002",
  "USGS:02291597:00011:00001",
  "USGS:02317620:00011:00001",
  "USGS:02317620:00011:00002",
  "USGS:02319000:00011:00002",
  "USGS:02319000:00011:00003",
  "USGS:02319300:00011:00004",
  "USGS:02319300:00011:00001",
  "USGS:02319302:00011:00016",
  "USGS:02319302:00011:00003",
  "USGS:02319302:00011:00002",
  "USGS:02319302:00011:00017",
  "USGS:02319302:00011:00018",
  "USGS:02319302:00011:00019",
  "USGS:02319302:00011:00020",
  "USGS:02319394:00011:00005",
  "USGS:02319394:00011:00004",
  "USGS:02319500:00011:00003",
  "USGS:02299472:00011:00012",
  "USGS:02299472:00011:00001",
  "USGS:02299472:00011:00002",
  "USGS:02299482:00011:00002",
  "USGS:02299482:00011:00005",
  "USGS:02299482:00011:00001",
  "USGS:02299482:00011:00004",
  "USGS:02299484:00011:00002",
  "USGS:02299484:00011:00001",
  "USGS:02299710:00011:00002",
  "USGS:02299710:00011:00001",
  "USGS:02299710:00011:00003",
  "USGS:02299710:00011:00004",
  "USGS:02299710:00011:00005",
  "USGS:02299727:00011:00003",
  "USGS:02299727:00011:00005",
  "USGS:02299727:00011:00001",
  "USGS:02299727:00011:00002",
  "USGS:02299727:00011:00004",
  "USGS:02299733:00011:00003",
  "USGS:02299733:00011:00005",
  "USGS:02299733:00011:00001",
  "USGS:02299733:00011:00002",
  "USGS:02299733:00011:00004",
  "USGS:02299735:00011:00003",
  "USGS:02299735:00011:00005",
  "USGS:02299735:00011:00001",
  "USGS:02299735:00011:00002",
  "USGS:02299735:00011:00004",
  "USGS:02299861:00011:00002",
  "USGS:02299861:00011:00001",
  "USGS:02299950:00011:00005",
  "USGS:02299950:00011:00002",
  "USGS:02299950:00011:00015",
  "USGS:023000095:00011:00013",
  "USGS:023000095:00011:00015",
  "USGS:023000095:00011:00002",
  "USGS:023000095:00011:00014",
  "USGS:023000095:00011:00016",
  "USGS:02300017:00011:00002",
  "USGS:02300017:00011:00001",
  "USGS:02300018:00011:00002",
  "USGS:02300018:00011:00001",
  "USGS:02300021:00011:00004",
  "USGS:02300021:00011:00005",
  "USGS:02300021:00011:00015",
  "USGS:02300021:00011:00023",
  "USGS:02300021:00011:00001",
  "USGS:02300021:00011:00002",
  "USGS:02300021:00011:00003",
  "USGS:02300021:00011:00026",
  "USGS:02300033:00011:00012",
  "USGS:02300033:00011:00011",
  "USGS:02300033:00011:00001",
  "USGS:02300042:00011:00002",
  "USGS:02300042:00011:00014",
  "USGS:02300042:00011:00013",
  "USGS:02300075:00011:00002",
  "USGS:02300075:00011:00001",
  "USGS:02300082:00011:00002",
  "USGS:02300082:00011:00004",
  "USGS:02300082:00011:00001",
  "USGS:02300100:00011:00001",
  "USGS:02300100:00011:00002",
  "USGS:02300100:00011:00012",
  "USGS:02300210:00011:00002",
  "USGS:02300210:00011:00001",
  "USGS:02300300:00011:00002",
  "USGS:02300300:00011:00001",
  "USGS:02300300:00011:00012",
  "USGS:02300500:00011:00007",
  "USGS:02300500:00011:00002",
  "USGS:02300500:00011:00003",
  "USGS:02300500:00011:00024",
  "USGS:02300700:00011:00001",
  "USGS:02300700:00011:00002",
  "USGS:02300700:00011:00015",
  "USGS:02300703:00011:00001",
  "USGS:02300882:00011:00002",
  "USGS:02300882:00011:00001",
  "USGS:02300995:00011:00001",
  "USGS:02301000:00011:00002",
  "USGS:02301000:00011:00003",
  "USGS:02301000:00011:00017",
  "USGS:02301150:00011:00012",
  "USGS:02301150:00011:00002",
  "USGS:02301150:00011:00001",
  "USGS:02301300:00011:00002",
  "USGS:02301300:00011:00003",
  "USGS:02301300:00011:00017",
  "USGS:02301500:00011:00004",
  "USGS:02301500:00011:00002",
  "USGS:02301500:00011:00003",
  "USGS:02301500:00011:00023",
  "USGS:02301638:00011:00002",
  "USGS:02301638:00011:00004",
  "USGS:02301638:00011:00001",
  "USGS:02301638:00011:00003",
  "USGS:02301638:00011:00005",
  "USGS:02301718:00011:00003",
  "USGS:02301718:00011:00005",
  "USGS:02301718:00011:00002",
  "USGS:02301718:00011:00004",
  "USGS:02301718:00011:00006",
  "USGS:02301719:00011:00003",
  "USGS:02301719:00011:00002",
  "USGS:02301719:00011:00005",
  "USGS:02301719:00011:00001",
  "USGS:02301719:00011:00004",
  "USGS:02301719:00011:00023",
  "USGS:02301721:00011:00006",
  "USGS:02301721:00011:00008",
  "USGS:02301721:00011:00031",
  "USGS:02301721:00011:00003",
  "USGS:02301721:00011:00007",
  "USGS:02301721:00011:00009",
  "USGS:02301721:00011:00030",
  "USGS:02301721:00011:00032",
  "USGS:02301738:00011:00002",
  "USGS:02301738:00011:00001",
  "USGS:02301740:00011:00002",
  "USGS:02301740:00011:00012",
  "USGS:02301740:00011:00001",
  "USGS:02301745:00011:00002",
  "USGS:02301745:00011:00012",
  "USGS:02301745:00011:00001",
  "USGS:02301750:00011:00003",
  "USGS:02301750:00011:00001",
  "USGS:02301750:00011:00002",
  "USGS:02301750:00011:00014",
  "USGS:02301793:00011:00002",
  "USGS:02301793:00011:00001",
  "USGS:02301900:00011:00001",
  "USGS:02301900:00011:00002",
  "USGS:02301990:00011:00001",
  "USGS:02301990:00011:00002",
  "USGS:02301990:00011:00013",
  "USGS:02302000:00011:00001",
  "USGS:02302000:00011:00013",
  "USGS:02302010:00011:00001",
  "USGS:02302010:00011:00002",
  "USGS:02302010:00011:00013",
  "USGS:02302500:00011:00013",
  "USGS:02302500:00011:00001",
  "USGS:02302500:00011:00002",
  "USGS:02303000:00011:00002",
  "USGS:02303000:00011:00003",
  "USGS:02303000:00011:00006",
  "USGS:02303205:00011:00002",
  "USGS:02303205:00011:00001",
  "USGS:02303330:00011:00014",
  "USGS:02303330:00011:00001",
  "USGS:02303330:00011:00002",
  "USGS:02303348:00011:00011",
  "USGS:02303348:00011:00001",
  "USGS:02357700:00011:00001",
  "USGS:02358000:00011:00026",
  "USGS:02358000:00011:00002",
  "USGS:02358000:00011:00003",
  "USGS:02358000:00011:00013",
  "USGS:02358700:00011:00001",
  "USGS:02358700:00011:00002",
  "USGS:02358789:00011:00003",
  "USGS:02358789:00011:00001",
  "USGS:02359000:00011:00010",
  "USGS:02359000:00011:00002",
  "USGS:02359000:00011:00003",
  "USGS:02359170:00011:00001",
  "USGS:02359170:00011:00002",
  "USGS:02359315:00011:00002",
  "USGS:02359315:00011:00001",
  "USGS:02359500:00011:00002",
  "USGS:02359500:00011:00003",
  "USGS:02365200:00011:00001",
  "USGS:02365200:00011:00002",
  "USGS:02365470:00011:00002",
  "USGS:02365470:00011:00001",
  "USGS:02303350:00011:00001",
  "USGS:02303350:00011:00002",
  "USGS:02303350:00011:00012",
  "USGS:02303400:00011:00002",
  "USGS:02303400:00011:00003",
  "USGS:02303400:00011:00014",
  "USGS:02303410:00011:00011",
  "USGS:02303410:00011:00001",
  "USGS:02303420:00011:00001",
  "USGS:02303420:00011:00002",
  "USGS:02303420:00011:00013",
  "USGS:02303424:00011:00001",
  "USGS:02303800:00011:00001",
  "USGS:02303800:00011:00002",
  "USGS:02304000:00011:00003",
  "USGS:02304000:00011:00002",
  "USGS:02304000:00011:00004",
  "USGS:02304000:00011:00005",
  "USGS:02304000:00011:00015",
  "USGS:02304500:00011:00009",
  "USGS:02304500:00011:00036",
  "USGS:02304500:00011:00002",
  "USGS:02304510:00011:00008",
  "USGS:02304510:00011:00009",
  "USGS:02304510:00011:00002",
  "USGS:02304510:00011:00006",
  "USGS:02304510:00011:00007",
  "USGS:02304510:00011:00018",
  "USGS:02304520:00011:00001",
  "USGS:02304520:00011:00003",
  "USGS:02304520:00011:00005",
  "USGS:02304520:00011:00007",
  "USGS:02304520:00011:00002",
  "USGS:02304520:00011:00004",
  "USGS:02304520:00011:00006",
  "USGS:02305851:00011:00002",
  "USGS:02305851:00011:00001",
  "USGS:02306000:00011:00013",
  "USGS:02306000:00011:00001",
  "USGS:02306000:00011:00002",
  "USGS:02306000:00011:00014",
  "USGS:02306000:00011:00016",
  "USGS:023060003:00011:00002",
  "USGS:023060003:00011:00012",
  "USGS:023060003:00011:00001",
  "USGS:023060003:00011:00003",
  "USGS:023060003:00011:00026",
  "USGS:02306028:00011:00012",
  "USGS:02306028:00011:00013",
  "USGS:02306028:00011:00015",
  "USGS:02306028:00011:00005",
  "USGS:02306028:00011:00009",
  "USGS:02306028:00011:00011",
  "USGS:02306028:00011:00014",
  "USGS:02306647:00011:00001",
  "USGS:02306647:00011:00002",
  "USGS:02306647:00011:00014",
  "USGS:02306654:00011:00001",
  "USGS:02306654:00011:00002",
  "USGS:02306774:00011:00001",
  "USGS:02306774:00011:00002",
  "USGS:02306774:00011:00014",
  "USGS:02306904:00011:00001",
  "USGS:02306950:00011:00003",
  "USGS:02306950:00011:00001",
  "USGS:02307032:00011:00002",
  "USGS:02307032:00011:00001",
  "USGS:02307032:00011:00013",
  "USGS:02307200:00011:00002",
  "USGS:02307200:00011:00003",
  "USGS:02307323:00011:00001",
  "USGS:02307323:00011:00002",
  "USGS:02307359:00011:00001",
  "USGS:02307359:00011:00002",
  "USGS:02307362:00011:00001",
  "USGS:02307445:00011:00002",
  "USGS:02307445:00011:00001",
  "USGS:02307498:00011:00019",
  "USGS:02307498:00011:00007",
  "USGS:02307498:00011:00008",
  "USGS:02307498:00011:00003",
  "USGS:02307498:00011:00004",
  "USGS:02307498:00011:00005",
  "USGS:02307498:00011:00006",
  "USGS:02307668:00011:00002",
  "USGS:02307668:00011:00001",
  "USGS:02307669:00011:00003",
  "USGS:02307669:00011:00001",
  "USGS:02307674:00011:00003",
  "USGS:02307674:00011:00002",
  "USGS:02307674:00011:00001",
  "USGS:02307780:00011:00001",
  "USGS:02307780:00011:00002",
  "USGS:02307834:00011:00002",
  "USGS:02307834:00011:00001",
  "USGS:02307835:00011:00001",
  "USGS:02307836:00011:00001",
  "USGS:02308861:00011:00001",
  "USGS:02308865:00011:00011",
  "USGS:02308865:00011:00001",
  "USGS:02308866:00011:00001",
  "USGS:02308870:00011:00003",
  "USGS:02308870:00011:00002",
  "USGS:02308870:00011:00001",
  "USGS:02308889:00011:00002",
  "USGS:02308935:00011:00001",
  "USGS:02308935:00011:00002",
  "USGS:02308935:00011:00003",
  "USGS:02309110:00011:00003",
  "USGS:02309110:00011:00002",
  "USGS:02309415:00011:00003",
  "USGS:02309415:00011:00002",
  "USGS:02309415:00011:00001",
  "USGS:02309421:00011:00002",
  "USGS:02309421:00011:00001",
  "USGS:02309425:00011:00003",
  "USGS:02309425:00011:00002",
  "USGS:02309425:00011:00001",
  "USGS:02309740:00011:00001",
  "USGS:02309848:00011:00001",
  "USGS:02309848:00011:00002",
  "USGS:02310000:00011:00002",
  "USGS:02310000:00011:00003",
  "USGS:02310075:00011:00001",
  "USGS:02310280:00011:00001",
  "USGS:02310280:00011:00002",
  "USGS:02310280:00011:00013",
  "USGS:02310286:00011:00002",
  "USGS:02310286:00011:00001",
  "USGS:02313231:00011:00002",
  "USGS:252612080300701:00011:00001",
  "USGS:252619080310201:00011:00001",
  "USGS:252718080264901:00011:00010",
  "USGS:252820080505401:00011:00003",
  "USGS:252820080505401:00011:00002",
  "USGS:252820080505401:00011:00004",
  "USGS:252820080505401:00011:00001",
  "USGS:252906080213101:00011:00001",
  "USGS:252918080234201:00011:00001",
  "USGS:252928080332401:00011:00001",
  "USGS:252933080210001:00011:00001",
  "USGS:253029080295601:00011:00002",
  "USGS:253044080555900:00011:00002",
  "USGS:253044080555900:00011:00001",
  "USGS:253044080555900:00011:00003",
  "USGS:253828080391100:00011:00003",
  "USGS:02236125:00011:00011",
  "USGS:02236160:00011:00004",
  "USGS:02236160:00011:00001",
  "USGS:02236160:00011:00011",
  "USGS:02236350:00011:00002",
  "USGS:02236350:00011:00003",
  "USGS:02236500:00011:00002",
  "USGS:02236500:00011:00003",
  "USGS:02236500:00011:00013",
  "USGS:02236605:00011:00001",
  "USGS:02236605:00011:00002",
  "USGS:02236840:00011:00001",
  "USGS:02236900:00011:00001",
  "USGS:02236900:00011:00002",
  "USGS:02236900:00011:00013",
  "USGS:02236900:00011:00014",
  "USGS:02236901:00011:00001",
  "USGS:02237000:00011:00001",
  "USGS:02237000:00011:00003",
  "USGS:02237001:00011:00001",
  "USGS:02237010:00011:00001",
  "USGS:02237011:00011:00001",
  "USGS:02237050:00011:00001",
  "USGS:02237051:00011:00001",
  "USGS:02237206:00011:00001",
  "USGS:02237207:00011:00001",
  "USGS:02237293:00011:00001",
  "USGS:02237293:00011:00002",
  "USGS:02237293:00011:00003",
  "USGS:02237698:00011:00003",
  "USGS:02237698:00011:00002",
  "USGS:02237698:00011:00001",
  "USGS:02237700:00011:00014",
  "USGS:02237700:00011:00012",
  "USGS:02237700:00011:00018",
  "USGS:02237700:00011:00002",
  "USGS:02237700:00011:00013",
  "USGS:02237700:00011:00008",
  "USGS:02237700:00011:00009",
  "USGS:02237700:00011:00020",
  "USGS:02237701:00011:00001",
  "USGS:02237701:00011:00002",
  "USGS:02237734:00011:00002",
  "USGS:02237734:00011:00001",
  "USGS:02238000:00011:00002",
  "USGS:02238000:00011:00003",
  "USGS:02238000:00011:00004",
  "USGS:02238000:00011:00010",
  "USGS:02238000:00011:00011",
  "USGS:02238000:00011:00012",
  "USGS:02238000:00011:00013",
  "USGS:02238000:00011:00016",
  "USGS:02238001:00011:00001",
  "USGS:02238001:00011:00002",
  "USGS:02238499:00011:00001",
  "USGS:02238499:00011:00002",
  "USGS:02238500:00011:00016",
  "USGS:02238500:00011:00003",
  "USGS:02238500:00011:00007",
  "USGS:02238500:00011:00008",
  "USGS:02238500:00011:00011",
  "USGS:02238500:00011:00012",
  "USGS:02238500:00011:00015",
  "USGS:02238500:00011:00019",
  "USGS:02239000:00011:00001",
  "USGS:02239000:00011:00002",
  "USGS:02239500:00011:00003",
  "USGS:02239500:00011:00010",
  "USGS:02239501:00011:00002",
  "USGS:02239501:00011:00001",
  "USGS:02239600:00011:00003",
  "USGS:02239600:00011:00001",
  "USGS:02239601:00011:00001",
  "USGS:02240000:00011:00002",
  "USGS:02240000:00011:00003",
  "USGS:02240000:00011:00008",
  "USGS:02240500:00011:00002",
  "USGS:02240500:00011:00003",
  "USGS:02240500:00011:00007",
  "USGS:02243000:00011:00002",
  "USGS:02243000:00011:00003",
  "USGS:02243000:00011:00005",
  "USGS:02243959:00011:00001",
  "USGS:02243959:00011:00002",
  "USGS:02243960:00011:00001",
  "USGS:02243960:00011:00002",
  "USGS:02243960:00011:00004",
  "USGS:02243960:00011:00005",
  "USGS:02243960:00011:00006",
  "USGS:02243960:00011:00007",
  "USGS:02243960:00011:00008",
  "USGS:02244040:00011:00016",
  "USGS:02244040:00011:00018",
  "USGS:02244040:00011:00001",
  "USGS:02244040:00011:00017",
  "USGS:02244040:00011:00015",
  "USGS:02244040:00011:00023",
  "USGS:02244333:00011:00002",
  "USGS:02244333:00011:00001",
  "USGS:02244440:00011:00001",
  "USGS:02244440:00011:00002",
  "USGS:02244440:00011:00012",
  "USGS:02245260:00011:00016",
  "USGS:02245260:00011:00005",
  "USGS:02245260:00011:00001",
  "USGS:02245260:00011:00017",
  "USGS:02245260:00011:00018",
  "USGS:02245260:00011:00009",
  "USGS:02245260:00011:00019",
  "USGS:02245500:00011:00001",
  "USGS:02245500:00011:00002",
  "USGS:02245500:00011:00004",
  "USGS:02246000:00011:00001",
  "USGS:02246000:00011:00002",
  "USGS:02246000:00011:00009",
  "USGS:02246010:00011:00002",
  "USGS:02246010:00011:00001",
  "USGS:02246500:00011:00002",
  "USGS:02246500:00011:00006",
  "USGS:02246500:00011:00022",
  "USGS:02247510:00011:00003",
  "USGS:02247510:00011:00004",
  "USGS:02247510:00011:00006",
  "USGS:02248000:00011:00002",
  "USGS:02248000:00011:00003",
  "USGS:02248000:00011:00005",
  "USGS:02248350:00011:00001",
  "USGS:02248350:00011:00008",
  "USGS:02248380:00011:00021",
  "USGS:02248380:00011:00003",
  "USGS:02248380:00011:00001",
  "USGS:02248380:00011:00022",
  "USGS:02248380:00011:00009",
  "USGS:02248380:00011:00012",
  "USGS:02248650:00011:00003",
  "USGS:02248650:00011:00001",
  "USGS:02248660:00011:00003",
  "USGS:02248660:00011:00001",
  "USGS:02249007:00011:00002",
  "USGS:02249007:00011:00001",
  "USGS:02249007:00011:00003",
  "USGS:254344081095101:00011:00003",
  "USGS:254344081095101:00011:00002",
  "USGS:254344081095101:00011:00004",
  "USGS:254344081095101:00011:00001",
  "USGS:254442080305201:00011:00001",
  "USGS:254445080295001:00011:00001",
  "USGS:254446080295501:00011:00001",
  "USGS:254543080405401:00011:00036",
  "USGS:254543080405401:00011:00024",
  "USGS:254543080405401:00011:00023",
  "USGS:254543080405401:00011:00031",
  "USGS:254543080405401:00011:00035",
  "USGS:254543080405401:00011:00048",
  "USGS:02310663:00011:00021",
  "USGS:02310663:00011:00002",
  "USGS:02310663:00011:00012",
  "USGS:02310663:00011:00025",
  "USGS:02310673:00011:00003",
  "USGS:02310673:00011:00005",
  "USGS:02310673:00011:00001",
  "USGS:02310673:00011:00002",
  "USGS:02310673:00011:00004",
  "USGS:02310674:00011:00003",
  "USGS:02310674:00011:00005",
  "USGS:02310674:00011:00001",
  "USGS:02310674:00011:00002",
  "USGS:02310674:00011:00004",
  "USGS:02310675:00011:00002",
  "USGS:02310678:00011:00024",
  "USGS:02310678:00011:00023",
  "USGS:02310678:00011:00002",
  "USGS:02310678:00011:00026",
  "USGS:02310678:00011:00025",
  "USGS:02310688:00011:00016",
  "USGS:02310688:00011:00018",
  "USGS:02310688:00011:00019",
  "USGS:02310688:00011:00001",
  "USGS:02310688:00011:00015",
  "USGS:02310688:00011:00017",
  "USGS:02310689:00011:00003",
  "USGS:02310689:00011:00005",
  "USGS:02310689:00011:00004",
  "USGS:02310689:00011:00018",
  "USGS:02310689:00011:00001",
  "USGS:02310689:00011:00002",
  "USGS:02310700:00011:00016",
  "USGS:02310700:00011:00027",
  "USGS:02310700:00011:00021",
  "USGS:02310700:00011:00030",
  "USGS:02310700:00011:00003",
  "USGS:02310700:00011:00015",
  "USGS:02310700:00011:00026",
  "USGS:02310700:00011:00029",
  "USGS:02310742:00011:00003",
  "USGS:02310742:00011:00007",
  "USGS:02310742:00011:00001",
  "USGS:02310742:00011:00002",
  "USGS:02310742:00011:00006",
  "USGS:02310747:00011:00007",
  "USGS:02310747:00011:00009",
  "USGS:02310747:00011:00003",
  "USGS:02310747:00011:00001",
  "USGS:02310747:00011:00008",
  "USGS:02310747:00011:00021",
  "USGS:02310752:00011:00003",
  "USGS:02310752:00011:00005",
  "USGS:02310752:00011:00001",
  "USGS:02310752:00011:00002",
  "USGS:02310752:00011:00004",
  "USGS:02310947:00011:00002",
  "USGS:02310947:00011:00003",
  "USGS:02311000:00011:00001",
  "USGS:02311000:00011:00002",
  "USGS:02311500:00011:00002",
  "USGS:02311500:00011:00003",
  "USGS:02312000:00011:00001",
  "USGS:02312000:00011:00002",
  "USGS:02312180:00011:00002",
  "USGS:02312180:00011:00003",
  "USGS:02312180:00011:00011",
  "USGS:02312200:00011:00002",
  "USGS:02312200:00011:00003",
  "USGS:02312300:00011:00013",
  "USGS:02312300:00011:00001",
  "USGS:02312500:00011:00001",
  "USGS:02312500:00011:00002",
  "USGS:02312558:00011:00013",
  "USGS:02312558:00011:00001",
  "USGS:02312598:00011:00001",
  "USGS:02312598:00011:00002",
  "USGS:02312600:00011:00001",
  "USGS:02312600:00011:00002",
  "USGS:02312640:00011:00002",
  "USGS:02312640:00011:00001",
  "USGS:02312645:00011:00001",
  "USGS:02312645:00011:00002",
  "USGS:02312667:00011:00001",
  "USGS:02312667:00011:00002",
  "USGS:02312667:00011:00005",
  "USGS:02312675:00011:00008",
  "USGS:02312675:00011:00001",
  "USGS:02312675:00011:00010",
  "USGS:02312700:00011:00001",
  "USGS:02312700:00011:00003",
  "USGS:02312700:00011:00019",
  "USGS:02312719:00011:00001",
  "USGS:02312719:00011:00003",
  "USGS:02312720:00011:00001",
  "USGS:02312720:00011:00002",
  "USGS:02312720:00011:00007",
  "USGS:02312722:00011:00001",
  "USGS:02312722:00011:00002",
  "USGS:02312722:00011:00004",
  "USGS:02312762:00011:00001",
  "USGS:02312762:00011:00002",
  "USGS:02312762:00011:00005",
  "USGS:02312764:00011:00004",
  "USGS:02312764:00011:00001",
  "USGS:02313000:00011:00002",
  "USGS:02313000:00011:00003",
  "USGS:02313000:00011:00013",
  "USGS:02313098:00011:00001",
  "USGS:02313100:00011:00012",
  "USGS:02313100:00011:00002",
  "USGS:02313100:00011:00003",
  "USGS:02313100:00011:00009",
  "USGS:02313200:00011:00002",
  "USGS:02313200:00011:00010",
  "USGS:02313230:00011:00002",
  "USGS:02313230:00011:00003",
  "USGS:02313230:00011:00005",
  "USGS:02313230:00011:00006",
  "USGS:02313250:00011:00002",
  "USGS:02313250:00011:00003",
  "USGS:02313250:00011:00005",
  "USGS:02313250:00011:00006",
  "USGS:02313272:00011:00006",
  "USGS:02313272:00011:00008",
  "USGS:02313272:00011:00004",
  "USGS:02313272:00011:00005",
  "USGS:02313272:00011:00007",
  "USGS:02313700:00011:00003",
  "USGS:02313700:00011:00004",
  "USGS:02315000:00011:00001",
  "USGS:02315000:00011:00002",
  "USGS:02315500:00011:00001",
  "USGS:02315500:00011:00002",
  "USGS:02315550:00011:00002",
  "USGS:02315550:00011:00001",
  "USGS:02315626:00011:00004",
  "USGS:02315626:00011:00001",
  "USGS:260355080541401:00011:00001",
  "USGS:260405081414101:00011:00001",
  "USGS:260410080452701:00011:00001",
  "USGS:260458080134801:00011:00001",
  "USGS:260536080302501:00011:00001",
  "USGS:260725080451001:00011:00001",
  "USGS:260810080222001:00011:00001",
  "USGS:260821080185101:00011:00001",
  "USGS:261023080443001:00011:00001",
  "USGS:02228500:00011:00005",
  "USGS:02231000:00011:00002",
  "USGS:02231000:00011:00003",
  "USGS:02231000:00011:00015",
  "USGS:02231291:00011:00002",
  "USGS:02231291:00011:00001",
  "USGS:02231291:00011:00003",
  "USGS:02231291:00011:00012",
  "USGS:02231342:00011:00001",
  "USGS:02231342:00011:00002",
  "USGS:02231342:00011:00004",
  "USGS:02231396:00011:00002",
  "USGS:02231396:00011:00001",
  "USGS:02231396:00011:00005",
  "USGS:02231454:00011:00002",
  "USGS:02231454:00011:00001",
  "USGS:02231454:00011:00004",
  "USGS:02231600:00011:00002",
  "USGS:02231600:00011:00003",
  "USGS:02231600:00011:00006",
  "USGS:02232000:00011:00002",
  "USGS:02232000:00011:00003",
  "USGS:02232000:00011:00008",
  "USGS:02232155:00011:00002",
  "USGS:02232155:00011:00001",
  "USGS:02232200:00011:00001",
  "USGS:02232200:00011:00002",
  "USGS:02232200:00011:00004",
  "USGS:02232400:00011:00001",
  "USGS:02232400:00011:00002",
  "USGS:02232400:00011:00003",
  "USGS:02232400:00011:00004",
  "USGS:02232400:00011:00008",
  "USGS:02232500:00011:00002",
  "USGS:02232500:00011:00003",
  "USGS:02232500:00011:00009",
  "USGS:02233200:00011:00001",
  "USGS:02233200:00011:00002",
  "USGS:02233200:00011:00008",
  "USGS:02233475:00011:00002",
  "USGS:02233475:00011:00001",
  "USGS:02233484:00011:00001",
  "USGS:02233484:00011:00002",
  "USGS:02233484:00011:00004",
  "USGS:02233500:00011:00001",
  "USGS:02233500:00011:00002",
  "USGS:02233500:00011:00004",
  "USGS:02234000:00011:00006",
  "USGS:02234000:00011:00001",
  "USGS:02234000:00011:00002",
  "USGS:02234000:00011:00007",
  "USGS:02234000:00011:00008",
  "USGS:02234000:00011:00009",
  "USGS:02234324:00011:00001",
  "USGS:02234324:00011:00002",
  "USGS:02234324:00011:00004",
  "USGS:02234344:00011:00002",
  "USGS:02234344:00011:00001",
  "USGS:02234384:00011:00001",
  "USGS:02234384:00011:00002",
  "USGS:02234384:00011:00004",
  "USGS:02234400:00011:00001",
  "USGS:02234400:00011:00002",
  "USGS:02234400:00011:00005",
  "USGS:02234435:00011:00001",
  "USGS:02234435:00011:00002",
  "USGS:02234435:00011:00011",
  "USGS:02234500:00011:00018",
  "USGS:02234500:00011:00002",
  "USGS:02234500:00011:00001",
  "USGS:02234500:00011:00017",
  "USGS:02234500:00011:00008",
  "USGS:02234500:00011:00009",
  "USGS:02234990:00011:00001",
  "USGS:02234990:00011:00002",
  "USGS:02234990:00011:00005",
  "USGS:02234990:00011:00004",
  "USGS:02235000:00011:00002",
  "USGS:02235000:00011:00003",
  "USGS:02235000:00011:00006",
  "USGS:02235200:00011:00001",
  "USGS:02235200:00011:00002",
  "USGS:02235200:00011:00005",
  "USGS:02235500:00011:00015",
  "USGS:02235500:00011:00017",
  "USGS:02235500:00011:00001",
  "USGS:02235500:00011:00016",
  "USGS:02235500:00011:00008",
  "USGS:02235500:00011:00057",
  "USGS:02235500:00011:00054",
  "USGS:02236000:00011:00004",
  "USGS:02236000:00011:00001",
  "USGS:02236000:00011:00002",
  "USGS:02236000:00011:00005",
  "USGS:02236000:00011:00007",
  "USGS:02236000:00011:00008",
  "USGS:431045078160401:00011:00001",
  "USGS:431227075233301:00011:00001",
  "USGS:431308078544501:00011:00001",
  "USGS:431359075235501:00011:00001",
  "USGS:431841074573201:00011:00001",
  "USGS:432148076225101:00011:00001",
  "USGS:432148076225102:00011:00001",
  "USGS:432832074122201:00011:00001",
  "USGS:433001073474701:00011:00001",
  "USGS:433112075091501:00011:00001",
  "USGS:433258073440201:00011:00001",
  "USGS:435253073440701:00011:00001",
  "USGS:440114075453701:00011:00001",
  "USGS:440939075191301:00011:00001",
  "USGS:441214075542101:00011:00001",
  "USGS:441644073315101:00011:00001",
  "USGS:444904074455201:00011:00001",
  "USGS:445052073350201:00011:00001",
  "USGS:445216074593001:00011:00001",
  "USGS:445511074103901:00011:00001",
  "USGS:445511074103902:00011:00001",
  "USGS:445805073380501:00011:00001",
  "USGS:262554081283801:00011:00001",
  "USGS:262605081425901:00011:00001",
  "USGS:262703081340201:00011:00001",
  "USGS:02319500:00011:00004",
  "USGS:02319800:00011:00002",
  "USGS:02319800:00011:00001",
  "USGS:02320000:00011:00001",
  "USGS:02320000:00011:00002",
  "USGS:02320250:00011:00011",
  "USGS:02320250:00011:00002",
  "USGS:02320250:00011:00012",
  "USGS:02320250:00011:00013",
  "USGS:02320250:00011:00014",
  "USGS:02320250:00011:00015",
  "USGS:02320500:00011:00002",
  "USGS:02320500:00011:00003",
  "USGS:02320700:00011:00001",
  "USGS:02320700:00011:00002",
  "USGS:02321000:00011:00001",
  "USGS:02321000:00011:00002",
  "USGS:02321500:00011:00002",
  "USGS:02321500:00011:00003",
  "USGS:02321898:00011:00012",
  "USGS:02321898:00011:00001",
  "USGS:02322500:00011:00001",
  "USGS:02322500:00011:00003",
  "USGS:02322688:00011:00014",
  "USGS:02322688:00011:00003",
  "USGS:02322688:00011:00002",
  "USGS:02322688:00011:00015",
  "USGS:02322688:00011:00017",
  "USGS:02322688:00011:00016",
  "USGS:02322688:00011:00019",
  "USGS:02322700:00011:00002",
  "USGS:02322700:00011:00001",
  "USGS:02322703:00011:00001",
  "USGS:02322800:00011:00003",
  "USGS:02322800:00011:00001",
  "USGS:02322800:00011:00025",
  "USGS:02323000:00011:00001",
  "USGS:02323000:00011:00002",
  "USGS:02323500:00011:00005",
  "USGS:02323500:00011:00007",
  "USGS:02323500:00011:00006",
  "USGS:02323502:00011:00020",
  "USGS:02323502:00011:00003",
  "USGS:02323502:00011:00002",
  "USGS:02323502:00011:00021",
  "USGS:02323502:00011:00022",
  "USGS:02323502:00011:00023",
  "USGS:02323502:00011:00024",
  "USGS:02323566:00011:00026",
  "USGS:02323566:00011:00002",
  "USGS:02323566:00011:00004",
  "USGS:02323566:00011:00003",
  "USGS:02323566:00011:00027",
  "USGS:02323566:00011:00028",
  "USGS:02323566:00011:00029",
  "USGS:02323566:00011:00030",
  "USGS:02323567:00011:00001",
  "USGS:02323590:00011:00001",
  "USGS:02323592:00011:00008",
  "USGS:02323592:00011:00010",
  "USGS:02323592:00011:00003",
  "USGS:02323592:00011:00002",
  "USGS:02323592:00011:00009",
  "USGS:02323592:00011:00011",
  "USGS:02323592:00011:00005",
  "USGS:02323592:00011:00006",
  "USGS:02324000:00011:00002",
  "USGS:02324000:00011:00003",
  "USGS:02324400:00011:00001",
  "USGS:02324400:00011:00002",
  "USGS:02324500:00011:00002",
  "USGS:02325000:00011:00001",
  "USGS:02325000:00011:00002",
  "USGS:02326000:00011:00001",
  "USGS:02326000:00011:00002",
  "USGS:02326500:00011:00001",
  "USGS:02326500:00011:00002",
  "USGS:02326526:00011:00002",
  "USGS:02326526:00011:00001",
  "USGS:02326550:00011:00003",
  "USGS:02326900:00011:00001",
  "USGS:02326900:00011:00002",
  "USGS:02326993:00011:00002",
  "USGS:02327022:00011:00002",
  "USGS:02327022:00011:00003",
  "USGS:02327022:00011:00001",
  "USGS:02327031:00011:00003",
  "USGS:02327031:00011:00010",
  "USGS:02327031:00011:00011",
  "USGS:02327031:00011:00028",
  "USGS:02327031:00011:00002",
  "USGS:02327031:00011:00004",
  "USGS:02327031:00011:00005",
  "USGS:02327033:00011:00002",
  "USGS:02327033:00011:00001",
  "USGS:02327100:00011:00003",
  "USGS:02327100:00011:00004",
  "USGS:02328522:00011:00002",
  "USGS:02328522:00011:00001",
  "USGS:02329000:00011:00002",
  "USGS:02329000:00011:00003",
  "USGS:02329500:00011:00001",
  "USGS:02329500:00011:00002",
  "USGS:02329600:00011:00001",
  "USGS:02329600:00011:00003",
  "USGS:02329900:00011:00005",
  "USGS:02330000:00011:00001",
  "USGS:02330000:00011:00002",
  "USGS:02330100:00011:00001",
  "USGS:02330100:00011:00002",
  "USGS:02330150:00011:00002",
  "USGS:02330150:00011:00001",
  "USGS:02330400:00011:00003",
  "USGS:02330400:00011:00001",
  "USGS:02357500:00011:00004",
  "USGS:02357500:00011:00003",
  "USGS:02357500:00011:00001",
  "USGS:07227420:00011:00001",
  "USGS:07227420:00011:00004",
  "USGS:07227420:00011:00002",
  "USGS:07227460:00011:00002",
  "USGS:07227460:00011:00001",
  "USGS:02293254:00011:00012",
  "USGS:02293254:00011:00014",
  "USGS:02293262:00011:00002",
  "USGS:02293262:00011:00001",
  "USGS:02293987:00011:00002",
  "USGS:02293987:00011:00001",
  "USGS:02294161:00011:00001",
  "USGS:02294161:00011:00002",
  "USGS:02294217:00011:00001",
  "USGS:02294217:00011:00002",
  "USGS:02294260:00011:00002",
  "USGS:02294260:00011:00001",
  "USGS:02294260:00011:00014",
  "USGS:02294290:00011:00016",
  "USGS:02294290:00011:00001",
  "USGS:02294290:00011:00002",
  "USGS:02294330:00011:00001",
  "USGS:02294330:00011:00002",
  "USGS:02294405:00011:00001",
  "USGS:02294405:00011:00002",
  "USGS:02294650:00011:00002",
  "USGS:02294650:00011:00003",
  "USGS:02294650:00011:00021",
  "USGS:02294898:00011:00002",
  "USGS:02294898:00011:00003",
  "USGS:02295163:00011:00002",
  "USGS:02295163:00011:00001",
  "USGS:02295194:00011:00001",
  "USGS:02295194:00011:00002",
  "USGS:02295420:00011:00001",
  "USGS:02295420:00011:00002",
  "USGS:02295520:00011:00001",
  "USGS:02295520:00011:00011",
  "USGS:02295580:00011:00012",
  "USGS:02295580:00011:00001",
  "USGS:02295580:00011:00011",
  "USGS:02295637:00011:00002",
  "USGS:02295637:00011:00003",
  "USGS:02296260:00011:00002",
  "USGS:02296260:00011:00001",
  "USGS:02296260:00011:00016",
  "USGS:02296500:00011:00001",
  "USGS:02296500:00011:00002",
  "USGS:02296750:00011:00002",
  "USGS:02296750:00011:00003",
  "USGS:02297100:00011:00014",
  "USGS:02297100:00011:00017",
  "USGS:02297100:00011:00001",
  "USGS:02297100:00011:00002",
  "USGS:02297100:00011:00015",
  "USGS:02297105:00011:00011",
  "USGS:02297105:00011:00001",
  "USGS:02297155:00011:00001",
  "USGS:02297155:00011:00002",
  "USGS:02297310:00011:00002",
  "USGS:02297310:00011:00003",
  "USGS:02297345:00011:00004",
  "USGS:02297345:00011:00005",
  "USGS:02297345:00011:00001",
  "USGS:02297345:00011:00002",
  "USGS:02297345:00011:00003",
  "USGS:02297350:00011:00002",
  "USGS:02297350:00011:00003",
  "USGS:02297350:00011:00001",
  "USGS:02297350:00011:00004",
  "USGS:02297350:00011:00005",
  "USGS:02297600:00011:00002",
  "USGS:02297600:00011:00001",
  "USGS:02297635:00011:00002",
  "USGS:02297635:00011:00022",
  "USGS:02297635:00011:00001",
  "USGS:02297635:00011:00003",
  "USGS:02298110:00011:00002",
  "USGS:02298110:00011:00001",
  "USGS:02298123:00011:00001",
  "USGS:02298123:00011:00016",
  "USGS:02298124:00011:00004",
  "USGS:02298124:00011:00005",
  "USGS:02298170:00011:00002",
  "USGS:02298170:00011:00021",
  "USGS:02298170:00011:00001",
  "USGS:02298170:00011:00003",
  "USGS:02298202:00011:00015",
  "USGS:02298202:00011:00001",
  "USGS:02298202:00011:00002",
  "USGS:02298202:00011:00014",
  "USGS:02298488:00011:00002",
  "USGS:02298488:00011:00001",
  "USGS:02298492:00011:00002",
  "USGS:02298492:00011:00001",
  "USGS:02298492:00011:00014",
  "USGS:02298494:00011:00001",
  "USGS:02298495:00011:00002",
  "USGS:02298495:00011:00001",
  "USGS:02298527:00011:00002",
  "USGS:02298527:00011:00001",
  "USGS:02298530:00011:00002",
  "USGS:02298530:00011:00001",
  "USGS:02298554:00011:00002",
  "USGS:02298554:00011:00001",
  "USGS:02298608:00011:00001",
  "USGS:02298608:00011:00002",
  "USGS:02298760:00011:00001",
  "USGS:02298760:00011:00002",
  "USGS:02298830:00011:00002",
  "USGS:02298830:00011:00003",
  "USGS:02298880:00011:00001",
  "USGS:02298880:00011:00002",
  "USGS:021720709:00011:00002",
  "USGS:021720709:00011:00001",
  "USGS:021720709:00011:00003",
  "USGS:021720709:00011:00004",
  "USGS:272020082194801:00011:00001",
  "USGS:272058082143701:00011:00001",
  "USGS:272127082323801:00011:00001",
  "USGS:272129082330202:00011:00001",
  "USGS:272356082181302:00011:00001",
  "USGS:272404082161701:00011:00001",
  "USGS:14145100:00011:00002",
  "USGS:02250030:00011:00001",
  "USGS:02250030:00011:00002",
  "USGS:02250030:00011:00011",
  "USGS:02250030:00011:00013",
  "USGS:02251000:00011:00002",
  "USGS:02251000:00011:00001",
  "USGS:02251000:00011:00006",
  "USGS:02251500:00011:00002",
  "USGS:02251500:00011:00001",
  "USGS:02251500:00011:00004",
  "USGS:02251767:00011:00002",
  "USGS:02251767:00011:00001",
  "USGS:02251767:00011:00004",
  "USGS:02251800:00011:00001",
  "USGS:02251800:00011:00002",
  "USGS:02252500:00011:00001",
  "USGS:02252500:00011:00002",
  "USGS:02252500:00011:00004",
  "USGS:02253000:00011:00002",
  "USGS:02253000:00011:00003",
  "USGS:02253000:00011:00009",
  "USGS:02253000:00011:00010",
  "USGS:02253500:00011:00002",
  "USGS:02253500:00011:00003",
  "USGS:02253500:00011:00001",
  "USGS:02255600:00011:00002",
  "USGS:02255600:00011:00001",
  "USGS:02256500:00011:00002",
  "USGS:02256500:00011:00003",
  "USGS:02257000:00011:00012",
  "USGS:02257000:00011:00001",
  "USGS:02262900:00011:00001",
  "USGS:02262900:00011:00002",
  "USGS:02263800:00011:00001",
  "USGS:02263800:00011:00002",
  "USGS:02263850:00011:00001",
  "USGS:02263868:00011:00001",
  "USGS:02263869:00011:00002",
  "USGS:02263869:00011:00001",
  "USGS:02263870:00011:00001",
  "USGS:02264000:00011:00003",
  "USGS:02264000:00011:00001",
  "USGS:02264000:00011:00002",
  "USGS:02264000:00011:00004",
  "USGS:02264000:00011:00005",
  "USGS:02264003:00011:00002",
  "USGS:02264003:00011:00001",
  "USGS:02264003:00011:00010",
  "USGS:02264003:00011:00011",
  "USGS:02264004:00011:00001",
  "USGS:02264030:00011:00002",
  "USGS:02264030:00011:00001",
  "USGS:02264051:00011:00002",
  "USGS:02264051:00011:00001",
  "USGS:02264060:00011:00003",
  "USGS:02264060:00011:00001",
  "USGS:02264061:00011:00001",
  "USGS:02264100:00011:00006",
  "USGS:02264100:00011:00001",
  "USGS:02264100:00011:00002",
  "USGS:02264100:00011:00007",
  "USGS:02264100:00011:00008",
  "USGS:02264141:00011:00001",
  "USGS:02264495:00011:00001",
  "USGS:02264495:00011:00002",
  "USGS:02266025:00011:00002",
  "USGS:02266025:00011:00001",
  "USGS:02266026:00011:00001",
  "USGS:02266200:00011:00003",
  "USGS:02266200:00011:00001",
  "USGS:02266200:00011:00002",
  "USGS:02266200:00011:00004",
  "USGS:02266200:00011:00005",
  "USGS:02266205:00011:00002",
  "USGS:02266205:00011:00001",
  "USGS:02266206:00011:00001",
  "USGS:02266291:00011:00002",
  "USGS:02266291:00011:00001",
  "USGS:02266291:00011:00005",
  "USGS:02266291:00011:00008",
  "USGS:02266292:00011:00001",
  "USGS:02266293:00011:00002",
  "USGS:02266293:00011:00001",
  "USGS:02266293:00011:00003",
  "USGS:02266294:00011:00001",
  "USGS:02266295:00011:00002",
  "USGS:02266295:00011:00001",
  "USGS:02266296:00011:00001",
  "USGS:02266300:00011:00001",
  "USGS:02266300:00011:00003",
  "USGS:02266300:00011:00004",
  "USGS:02266300:00011:00005",
  "USGS:02266300:00011:00006",
  "USGS:02266480:00011:00001",
  "USGS:02266480:00011:00002",
  "USGS:02266495:00011:00001",
  "USGS:02266495:00011:00004",
  "USGS:02266495:00011:00002",
  "USGS:02266495:00011:00003",
  "USGS:02266496:00011:00003",
  "USGS:02266496:00011:00001",
  "USGS:02266550:00011:00001",
  "USGS:02266650:00011:00001",
  "USGS:02268400:00011:00001",
  "USGS:02268600:00011:00001",
  "USGS:02269148:00011:00001",
  "USGS:02269600:00011:00001",
  "USGS:02270000:00011:00001",
  "USGS:02270000:00011:00002",
  "USGS:14091500:00011:00001",
  "USGS:14091500:00011:00002",
  "USGS:14091500:00011:00003",
  "USGS:14092050:00011:00001",
  "USGS:14092500:00011:00001",
  "USGS:14092500:00011:00002",
  "USGS:14092500:00011:00003",
  "USGS:14092750:00011:00001",
  "USGS:14092750:00011:00002",
  "USGS:14093000:00011:00001",
  "USGS:14093000:00011:00002",
  "USGS:14096850:00011:00001",
  "USGS:14096850:00011:00002",
  "USGS:14097100:00011:00001",
  "USGS:254543080405401:00011:00033",
  "USGS:254543080405401:00011:00034",
  "USGS:254543080405401:00011:00037",
  "USGS:254543080491101:00011:00015",
  "USGS:254543080491101:00011:00023",
  "USGS:254543080491101:00011:00006",
  "USGS:254543080491101:00011:00007",
  "USGS:254720080253002:00011:00001",
  "USGS:254752080181501:00011:00001",
  "USGS:254754080344300:00011:00001",
  "USGS:254754080344300:00011:00003",
  "USGS:254759080483201:00011:00001",
  "USGS:254823080163701:00011:00001",
  "USGS:254823080175201:00011:00001",
  "USGS:254830080284201:00011:00001",
  "USGS:254848080432001:00011:00001",
  "USGS:254943080121501:00011:00001",
  "USGS:255014080355801:00011:00001",
  "USGS:255026080231300:00011:00001",
  "USGS:255026080240302:00011:00001",
  "USGS:255027080245501:00011:00001",
  "USGS:255030080221401:00011:00001",
  "USGS:255035080255401:00011:00001",
  "USGS:255036080270501:00011:00001",
  "USGS:255154080371300:00011:00015",
  "USGS:255154080371300:00011:00018",
  "USGS:255154080371300:00011:00005",
  "USGS:255154080371300:00011:00010",
  "USGS:255154080371300:00011:00030",
  "USGS:255154080371300:00011:00001",
  "USGS:255154080371300:00011:00014",
  "USGS:255154080371300:00011:00017",
  "USGS:255154080371300:00011:00013",
  "USGS:255154080371300:00011:00016",
  "USGS:255154080371300:00011:00019",
  "USGS:255154080371300:00011:00020",
  "USGS:255154080371300:00011:00002",
  "USGS:255154080371300:00011:00011",
  "USGS:255154080371300:00011:00007",
  "USGS:255154080371300:00011:00012",
  "USGS:255200080405001:00011:00011",
  "USGS:255200080405001:00011:00001",
  "USGS:255200080405001:00011:00012",
  "USGS:255200080405001:00011:00013",
  "USGS:255208080274001:00011:00001",
  "USGS:255209080212801:00011:00002",
  "USGS:255250080335001:00011:00001",
  "USGS:255300080370001:00011:00016",
  "USGS:255300080370001:00011:00017",
  "USGS:255300080370001:00011:00001",
  "USGS:255300080370001:00011:00012",
  "USGS:255300080370001:00011:00018",
  "USGS:255300080370001:00011:00019",
  "USGS:255300080370001:00011:00020",
  "USGS:255300080370001:00011:00021",
  "USGS:255300080370001:00011:00014",
  "USGS:255300080370001:00011:00015",
  "USGS:255327081275900:00011:00013",
  "USGS:255327081275900:00011:00003",
  "USGS:255327081275900:00011:00005",
  "USGS:255327081275900:00011:00012",
  "USGS:255327081275900:00011:00014",
  "USGS:255327081275900:00011:00009",
  "USGS:255358080260901:00011:00001",
  "USGS:255432081303900:00011:00012",
  "USGS:255432081303900:00011:00003",
  "USGS:255432081303900:00011:00005",
  "USGS:255432081303900:00011:00001",
  "USGS:255432081303900:00011:00014",
  "USGS:255437080103201:00011:00001",
  "USGS:255526080143001:00011:00002",
  "USGS:255534081324000:00011:00015",
  "USGS:255534081324000:00011:00019",
  "USGS:255534081324000:00011:00005",
  "USGS:255534081324000:00011:00012",
  "USGS:255534081324000:00011:00017",
  "USGS:255616080180301:00011:00001",
  "USGS:255634080450001:00011:00001",
  "USGS:255654081350200:00011:00014",
  "USGS:255654081350200:00011:00003",
  "USGS:255654081350200:00011:00005",
  "USGS:255654081350200:00011:00019",
  "USGS:255654081350200:00011:00016",
  "USGS:255708080295501:00011:00001",
  "USGS:255709080223701:00011:00001",
  "USGS:255726081303700:00011:00003",
  "USGS:255726081303700:00011:00007",
  "USGS:255726081303700:00011:00012",
  "USGS:255726081303700:00011:00013",
  "USGS:255726081303700:00011:00014",
  "USGS:255726081303700:00011:00015",
  "USGS:255726081303700:00011:00016",
  "USGS:255726081303700:00011:00017",
  "USGS:255726081303700:00011:00018",
  "USGS:255726081303700:00011:00011",
  "USGS:255726081303700:00011:00008",
  "USGS:255726081303700:00011:00010",
  "USGS:255726081303700:00011:00002",
  "USGS:255726081303700:00011:00006",
  "USGS:255732081363700:00011:00008",
  "USGS:255732081363700:00011:00013",
  "USGS:255732081363700:00011:00012",
  "USGS:255732081363700:00011:00007",
  "USGS:255828080401301:00011:00001",
  "USGS:260007080464401:00011:00001",
  "USGS:260010080085001:00011:00002",
  "USGS:260037080303401:00011:00001",
  "USGS:260042080351701:00011:00001",
  "USGS:260053080105701:00011:00001",
  "USGS:260111081243901:00011:00001",
  "USGS:260309081272601:00011:00001",
  "USGS:07227500:00011:00021",
  "USGS:260325080113901:00011:00001",
  "USGS:14155500:00011:00003",
  "USGS:14155500:00011:00001",
  "USGS:14155500:00011:00002",
  "USGS:14157500:00011:00002",
  "USGS:14157500:00011:00003",
  "USGS:14158100:00011:00001",
  "USGS:14158100:00011:00004",
  "USGS:14158100:00011:00002",
  "USGS:14158500:00011:00001",
  "USGS:14158500:00011:00002",
  "USGS:14158790:00011:00001",
  "USGS:14158790:00011:00002",
  "USGS:14158850:00011:00002",
  "USGS:14158850:00011:00004",
  "USGS:14159200:00011:00001",
  "USGS:14159200:00011:00002",
  "USGS:14159200:00011:00003",
  "USGS:14159400:00011:00002",
  "USGS:14159410:00011:00001",
  "USGS:14159500:00011:00001",
  "USGS:14159500:00011:00015",
  "USGS:14159500:00011:00016",
  "USGS:14159500:00011:00002",
  "USGS:14159500:00011:00003",
  "USGS:14159500:00011:00013",
  "USGS:14161100:00011:00002",
  "USGS:14161100:00011:00003",
  "USGS:14161500:00011:00001",
  "USGS:272504081120101:00011:00002",
  "USGS:272524080221800:00011:00015",
  "USGS:272524080221800:00011:00021",
  "USGS:272524080221800:00011:00001",
  "USGS:272524080242801:00011:00001",
  "USGS:272655080401601:00011:00001",
  "USGS:272838082142201:00011:00001",
  "USGS:273109080270301:00011:00001",
  "USGS:273126082384700:00011:00003",
  "USGS:273126082384700:00011:00005",
  "USGS:273126082384700:00011:00001",
  "USGS:273126082384700:00011:00002",
  "USGS:273126082384700:00011:00004",
  "USGS:273718082315501:00011:00001",
  "USGS:274812081190301:00011:00002",
  "USGS:275021082450500:00011:00001",
  "USGS:275815082440401:00011:00012",
  "USGS:275815082440401:00011:00001",
  "USGS:275917082222500:00011:00001",
  "USGS:280353082283400:00011:00001",
  "USGS:280842082392000:00011:00001",
  "USGS:281202081391701:00011:00001",
  "USGS:281448082301801:00011:00002",
  "USGS:281558082264601:00011:00001",
  "USGS:281714081093001:00011:00002",
  "USGS:282202081384601:00011:00002",
  "USGS:282202081384602:00011:00002",
  "USGS:282341081040101:00011:00002",
  "USGS:282406081093602:00011:00002",
  "USGS:282406081093602:00011:00001",
  "USGS:282434081283102:00011:00001",
  "USGS:282528081340901:00011:00001",
  "USGS:282531081082202:00011:00001",
  "USGS:282531081095701:00011:00002",
  "USGS:282532081075601:00011:00002",
  "USGS:282623081153801:00011:00002",
  "USGS:282738081341401:00011:00001",
  "USGS:282835081305201:00011:00001",
  "USGS:283154082313701:00011:00002",
  "USGS:283154082313701:00011:00001",
  "USGS:283249081053201:00011:00002",
  "USGS:284254081021000:00011:00001",
  "USGS:284551082345301:00011:00001",
  "USGS:284759081232100:00011:00001",
  "USGS:285531082412600:00011:00003",
  "USGS:285531082412600:00011:00005",
  "USGS:285531082412600:00011:00007",
  "USGS:285531082412600:00011:00001",
  "USGS:285531082412600:00011:00002",
  "USGS:285531082412600:00011:00004",
  "USGS:285531082412600:00011:00006",
  "USGS:290514082270701:00011:00002",
  "USGS:291100082010003:00011:00002",
  "USGS:291830081362200:00011:00001",
  "USGS:291830081362200:00011:00002",
  "USGS:291830081362200:00011:00003",
  "USGS:291830081362200:00011:00010",
  "USGS:291830081362200:00011:00013",
  "USGS:291830081362200:00011:00011",
  "USGS:292921082583285:00011:00002",
  "USGS:294213081345300:00011:00012",
  "USGS:294213081345300:00011:00013",
  "USGS:294213081345300:00011:00014",
  "USGS:294213081345300:00011:00015",
  "USGS:294213081345300:00011:00017",
  "USGS:294213081345300:00011:00016",
  "USGS:300010082594201:00011:00001",
  "USGS:300740084293001:00011:00002",
  "USGS:14187000:00011:00001",
  "USGS:14187000:00011:00002",
  "USGS:14187200:00011:00001",
  "USGS:14187200:00011:00002",
  "USGS:14187200:00011:00003",
  "USGS:14187500:00011:00002",
  "USGS:14187500:00011:00003",
  "USGS:14187600:00011:00002",
  "USGS:14187600:00011:00001",
  "USGS:14188610:00011:00002",
  "USGS:14188610:00011:00001",
  "USGS:14188800:00011:00002",
  "USGS:14188800:00011:00003",
  "USGS:14189000:00011:00002",
  "USGS:14189000:00011:00003",
  "USGS:14189050:00011:00001",
  "USGS:261035080221701:00011:00001",
  "USGS:261117080315201:00011:00001",
  "USGS:261141080163401:00011:00001",
  "USGS:261150080270001:00011:00001",
  "USGS:261150080270001:00011:00002",
  "USGS:261150080270001:00011:00005",
  "USGS:261150080270001:00011:00016",
  "USGS:261200080275001:00011:00001",
  "USGS:261200080275001:00011:00002",
  "USGS:261200080275001:00011:00004",
  "USGS:261200080275001:00011:00013",
  "USGS:261300080280001:00011:00001",
  "USGS:261300080280001:00011:00002",
  "USGS:261300080280001:00011:00013",
  "USGS:261300080280001:00011:00014",
  "USGS:261319080353201:00011:00001",
  "USGS:261347081351201:00011:00001",
  "USGS:261347081351202:00011:00001",
  "USGS:261347081351701:00011:00001",
  "USGS:261501080060701:00011:00001",
  "USGS:261533080571600:00011:00011",
  "USGS:261533080571600:00011:00068",
  "USGS:261533080571600:00011:00022",
  "USGS:261533080571600:00011:00001",
  "USGS:261533080571600:00011:00084",
  "USGS:261533080571600:00011:00083",
  "USGS:261533080571600:00011:00085",
  "USGS:261533080571600:00011:00082",
  "USGS:261533080571600:00011:00057",
  "USGS:261534080165801:00011:00001",
  "USGS:261543080495000:00011:00012",
  "USGS:261543080495000:00011:00005",
  "USGS:261543080495000:00011:00001",
  "USGS:261620081464402:00011:00001",
  "USGS:261641080064801:00011:00001",
  "USGS:261710080190001:00011:00001",
  "USGS:261735080534001:00011:00001",
  "USGS:261735080534002:00011:00001",
  "USGS:261808081042800:00011:00002",
  "USGS:261808081042800:00011:00001",
  "USGS:261808081042800:00011:00013",
  "USGS:261831080151301:00011:00001",
  "USGS:261903080065601:00011:00002",
  "USGS:261938080101001:00011:00001",
  "USGS:261957081432201:00011:00001",
  "USGS:261957081432202:00011:00001",
  "USGS:262038080584600:00011:00003",
  "USGS:262038080584600:00011:00002",
  "USGS:262038080584600:00011:00001",
  "USGS:262038080584600:00011:00033",
  "USGS:262100080190001:00011:00001",
  "USGS:262100080190001:00011:00002",
  "USGS:262100080190001:00011:00004",
  "USGS:262100080190001:00011:00013",
  "USGS:262158081283401:00011:00001",
  "USGS:262158081283402:00011:00001",
  "USGS:262158081283403:00011:00001",
  "USGS:262158081283404:00011:00001",
  "USGS:262200080210001:00011:00001",
  "USGS:262200080210001:00011:00002",
  "USGS:262200080210001:00011:00004",
  "USGS:262200080210001:00011:00013",
  "USGS:262212081312501:00011:00001",
  "USGS:262228081361901:00011:00001",
  "USGS:262240080258001:00011:00001",
  "USGS:262248081314101:00011:00001",
  "USGS:262258080273501:00011:00001",
  "USGS:262258081471802:00011:00001",
  "USGS:262300080220001:00011:00001",
  "USGS:262300080220001:00011:00002",
  "USGS:262300080220001:00011:00015",
  "USGS:262300080220001:00011:00016",
  "USGS:262317080074601:00011:00001",
  "USGS:262528080202700:00011:00001",
  "USGS:14299800:00011:00003",
  "USGS:14299800:00011:00002",
  "USGS:14299800:00011:00001",
  "USGS:14301000:00011:00006",
  "USGS:14301000:00011:00002",
  "USGS:14301000:00011:00004",
  "USGS:14301500:00011:00008",
  "USGS:14301500:00011:00001",
  "USGS:14301500:00011:00002",
  "USGS:14301500:00011:00009",
  "USGS:14301500:00011:00013",
  "USGS:14097100:00011:00002",
  "USGS:14103000:00011:00001",
  "USGS:14103000:00011:00002",
  "USGS:14103000:00011:00005",
  "USGS:14105700:00011:00021",
  "USGS:14105700:00011:00022",
  "USGS:14105700:00011:00023",
  "USGS:14105700:00011:00005",
  "USGS:14105700:00011:00002",
  "USGS:14105700:00011:00004",
  "USGS:14105700:00011:00012",
  "USGS:14105700:00011:00025",
  "USGS:14105800:00011:00001",
  "USGS:14113200:00011:00001",
  "USGS:14113200:00011:00002",
  "USGS:14113290:00011:00001",
  "USGS:14120000:00011:00001",
  "USGS:14120000:00011:00003",
  "USGS:14128870:00011:00001",
  "USGS:14137000:00011:00001",
  "USGS:14137000:00011:00002",
  "USGS:14138560:00011:00001",
  "USGS:14138720:00011:00012",
  "USGS:14138720:00011:00002",
  "USGS:14138720:00011:00001",
  "USGS:14138720:00011:00013",
  "USGS:14138800:00011:00001",
  "USGS:14138800:00011:00003",
  "USGS:14138850:00011:00005",
  "USGS:14138850:00011:00006",
  "USGS:14138850:00011:00004",
  "USGS:14138850:00011:00007",
  "USGS:14138870:00011:00005",
  "USGS:14138870:00011:00006",
  "USGS:14138870:00011:00021",
  "USGS:14138870:00011:00007",
  "USGS:14138900:00011:00005",
  "USGS:14138900:00011:00006",
  "USGS:14138900:00011:00004",
  "USGS:14138900:00011:00007",
  "USGS:14139000:00011:00001",
  "USGS:14139800:00011:00006",
  "USGS:14139800:00011:00022",
  "USGS:14139900:00011:00001",
  "USGS:14140000:00011:00001",
  "USGS:14140000:00011:00002",
  "USGS:14140020:00011:00001",
  "USGS:14141500:00011:00004",
  "USGS:14141500:00011:00001",
  "USGS:14141500:00011:00002",
  "USGS:14142500:00011:00003",
  "USGS:14142500:00011:00001",
  "USGS:14142800:00011:00002",
  "USGS:14142800:00011:00001",
  "USGS:14144800:00011:00001",
  "USGS:14144800:00011:00004",
  "USGS:14144900:00011:00001",
  "USGS:14144900:00011:00004",
  "USGS:14145110:00011:00001",
  "USGS:14145500:00011:00001",
  "USGS:14145500:00011:00002",
  "USGS:14145500:00011:00003",
  "USGS:14147500:00011:00003",
  "USGS:14147500:00011:00002",
  "USGS:14147500:00011:00004",
  "USGS:14148000:00011:00001",
  "USGS:14148000:00011:00002",
  "USGS:14148000:00011:00004",
  "USGS:14149000:00011:00002",
  "USGS:14149010:00011:00001",
  "USGS:14149500:00011:00001",
  "USGS:14149510:00011:00001",
  "USGS:14150000:00011:00001",
  "USGS:14150000:00011:00002",
  "USGS:14150000:00011:00008",
  "USGS:14150290:00011:00003",
  "USGS:14150290:00011:00001",
  "USGS:14150800:00011:00001",
  "USGS:14150800:00011:00002",
  "USGS:14150800:00011:00003",
  "USGS:14150900:00011:00002",
  "USGS:14151000:00011:00001",
  "USGS:14151000:00011:00002",
  "USGS:14151000:00011:00003",
  "USGS:14151000:00011:00005",
  "USGS:14151000:00011:00006",
  "USGS:14152000:00011:00001",
  "USGS:14152000:00011:00002",
  "USGS:14152000:00011:00003",
  "USGS:14152000:00011:00008",
  "USGS:14152000:00011:00007",
  "USGS:14153000:00011:00002",
  "USGS:14153500:00011:00003",
  "USGS:14153500:00011:00001",
  "USGS:14153500:00011:00002",
  "USGS:14154500:00011:00001",
  "USGS:14154500:00011:00002",
  "USGS:14155000:00011:00002",
  "USGS:06356500:00011:00001",
  "USGS:06356500:00011:00007",
  "USGS:06357800:00011:00001",
  "USGS:06357800:00011:00006",
  "USGS:06357800:00011:00003",
  "USGS:06359500:00011:00008",
  "USGS:06359500:00011:00002",
  "USGS:06359500:00011:00012",
  "USGS:06360500:00011:00001",
  "USGS:06360500:00011:00006",
  "USGS:06360500:00011:00003",
  "USGS:06395000:00011:00002",
  "USGS:06395000:00011:00003",
  "USGS:06395000:00011:00004",
  "USGS:06400000:00011:00006",
  "USGS:06400000:00011:00002",
  "USGS:06400000:00011:00003",
  "USGS:06400875:00011:00009",
  "USGS:06400875:00011:00001",
  "USGS:253044080555900:00011:00015",
  "USGS:253047080555600:00011:00013",
  "USGS:253047080555600:00011:00019",
  "USGS:253047080555600:00011:00020",
  "USGS:253047080555600:00011:00026",
  "USGS:253047080555600:00011:00001",
  "USGS:253047080555600:00011:00014",
  "USGS:253047080555600:00011:00015",
  "USGS:253047080555600:00011:00037",
  "USGS:253400080340401:00011:00001",
  "USGS:253413080225301:00011:00008",
  "USGS:253413080225301:00011:00007",
  "USGS:253413080225302:00011:00001",
  "USGS:253417080224301:00011:00008",
  "USGS:253417080224301:00011:00007",
  "USGS:253417080224302:00011:00001",
  "USGS:253419080223701:00011:00001",
  "USGS:253537080284401:00011:00001",
  "USGS:253539080320501:00011:00003",
  "USGS:253539080320501:00011:00001",
  "USGS:253632080321101:00011:00011",
  "USGS:253632080321101:00011:00001",
  "USGS:253644081013001:00011:00003",
  "USGS:253644081013001:00011:00002",
  "USGS:253644081013001:00011:00004",
  "USGS:253644081013001:00011:00001",
  "USGS:253708080304201:00011:00011",
  "USGS:253708080304201:00011:00001",
  "USGS:253828080391100:00011:00001",
  "USGS:253902080202501:00011:00002",
  "USGS:253937080304001:00011:00003",
  "USGS:253937080304001:00011:00001",
  "USGS:253948080250701:00011:00001",
  "USGS:253952080321501:00011:00001",
  "USGS:254000080181002:00011:00001",
  "USGS:254000080460001:00011:00001",
  "USGS:254054080295401:00011:00001",
  "USGS:254111080272501:00011:00001",
  "USGS:254112080294201:00011:00001",
  "USGS:254130080234501:00011:00002",
  "USGS:254130080380500:00011:00001",
  "USGS:254130080380500:00011:00004",
  "USGS:254138080284401:00011:00001",
  "USGS:254152080274501:00011:00001",
  "USGS:254152080282101:00011:00001",
  "USGS:254152080282601:00011:00001",
  "USGS:254157080213800:00011:00015",
  "USGS:254157080213800:00011:00016",
  "USGS:254157080213800:00011:00009",
  "USGS:254157080213800:00011:00001",
  "USGS:254158080294501:00011:00001",
  "USGS:254206080294701:00011:00001",
  "USGS:254207080300201:00011:00001",
  "USGS:254210080304801:00011:00001",
  "USGS:254213080281501:00011:00001",
  "USGS:254215080201503:00011:00001",
  "USGS:254218080241801:00011:00001",
  "USGS:254315080331500:00011:00001",
  "USGS:254315080331500:00011:00003",
  "USGS:254334080284401:00011:00001",
  "USGS:254340080203601:00011:00001",
  "USGS:254707080370201:00011:00001",
  "USGS:05051500:00011:00018",
  "USGS:05051500:00011:00003",
  "USGS:06403700:00011:00004",
  "USGS:06403700:00011:00002",
  "USGS:06403700:00011:00001",
  "USGS:06404000:00011:00008",
  "USGS:06404000:00011:00001",
  "USGS:06404000:00011:00007",
  "USGS:06404998:00011:00006",
  "USGS:06404998:00011:00001",
  "USGS:06404998:00011:00004",
  "USGS:06406000:00011:00006",
  "USGS:06406000:00011:00001",
  "USGS:06406000:00011:00004",
  "USGS:06406500:00011:00006",
  "USGS:06406500:00011:00002",
  "USGS:06406500:00011:00004",
  "USGS:06407500:00011:00007",
  "USGS:06407500:00011:00002",
  "USGS:06407500:00011:00006",
  "USGS:06408650:00011:00003",
  "USGS:06408650:00011:00002",
  "USGS:06408650:00011:00001",
  "USGS:06408700:00011:00002",
  "USGS:06408700:00011:00007",
  "USGS:06409000:00011:00010",
  "USGS:07227500:00011:00009",
  "USGS:07227500:00011:00008",
  "USGS:07227500:00011:00007",
  "USGS:07227500:00011:00020",
  "USGS:07227890:00011:00003",
  "USGS:07227890:00011:00005",
  "USGS:07227890:00011:00001",
  "USGS:07227900:00011:00002",
  "USGS:07227900:00011:00001",
  "USGS:07228000:00011:00003",
  "USGS:07228000:00011:00001",
  "USGS:07228000:00011:00002",
  "USGS:07233500:00011:00004",
  "USGS:07233500:00011:00001",
  "USGS:07233500:00011:00003",
  "USGS:11507500:00011:00003",
  "USGS:11507500:00011:00001",
  "USGS:11507500:00011:00002",
  "USGS:11507501:00011:00002",
  "USGS:11507501:00011:00005",
  "USGS:11507501:00011:00006",
  "USGS:11507501:00011:00003",
  "USGS:11507501:00011:00004",
  "USGS:11509105:00011:00002",
  "USGS:11509105:00011:00003",
  "USGS:11509105:00011:00011",
  "USGS:11509200:00011:00001",
  "USGS:11509200:00011:00010",
  "USGS:11509200:00011:00013",
  "USGS:11509250:00011:00001",
  "USGS:11509250:00011:00005",
  "USGS:11509340:00011:00007",
  "USGS:11509340:00011:00009",
  "USGS:11509340:00011:00001",
  "USGS:11509370:00011:00001",
  "USGS:11509370:00011:00004",
  "USGS:11509370:00011:00005",
  "USGS:11509370:00011:00002",
  "USGS:11509370:00011:00003",
  "USGS:11509500:00011:00012",
  "USGS:11509500:00011:00001",
  "USGS:11509500:00011:00002",
  "USGS:11510700:00011:00001",
  "USGS:11510700:00011:00002",
  "USGS:13181000:00011:00001",
  "USGS:13181000:00011:00002",
  "USGS:13183000:00011:00002",
  "USGS:13183000:00011:00001",
  "USGS:13215000:00011:00002",
  "USGS:13215000:00011:00001",
  "USGS:13217500:00011:00002",
  "USGS:13217500:00011:00001",
  "USGS:13233300:00011:00002",
  "USGS:13233300:00011:00001",
  "USGS:13290450:00011:00014",
  "USGS:13290450:00011:00015",
  "USGS:13331500:00011:00001",
  "USGS:13331500:00011:00002",
  "USGS:13331500:00011:00003",
  "USGS:13333000:00011:00001",
  "USGS:13333000:00011:00006",
  "USGS:14020000:00011:00002",
  "USGS:14020000:00011:00003",
  "USGS:14020300:00011:00001",
  "USGS:14020300:00011:00002",
  "USGS:14020850:00011:00001",
  "USGS:14020850:00011:00002",
  "USGS:14033500:00011:00002",
  "USGS:14033500:00011:00005",
  "USGS:14034470:00011:00006",
  "USGS:14034470:00011:00001",
  "USGS:14034470:00011:00002",
  "USGS:14034490:00011:00001",
  "USGS:14034500:00011:00001",
  "USGS:14034500:00011:00002",
  "USGS:14034500:00011:00005",
  "USGS:14034608:00011:00001",
  "USGS:14034608:00011:00002",
  "USGS:14036860:00011:00001",
  "USGS:14036860:00011:00002",
  "USGS:14038530:00011:00001",
  "USGS:14038530:00011:00002",
  "USGS:14043840:00011:00002",
  "USGS:14043840:00011:00001",
  "USGS:14044000:00011:00002",
  "USGS:14044000:00011:00003",
  "USGS:14046000:00011:00002",
  "USGS:14046000:00011:00003",
  "USGS:14046500:00011:00005",
  "USGS:14046500:00011:00006",
  "USGS:14046778:00011:00003",
  "USGS:14046778:00011:00002",
  "USGS:14046778:00011:00001",
  "USGS:14046890:00011:00003",
  "USGS:14046890:00011:00004",
  "USGS:14046890:00011:00002",
  "USGS:14046890:00011:00001",
  "USGS:14048000:00011:00002",
  "USGS:14048000:00011:00008",
  "USGS:14076500:00011:00001",
  "USGS:14076500:00011:00002",
  "USGS:14076500:00011:00003",
  "USGS:14087380:00011:00003",
  "USGS:14087380:00011:00002",
  "USGS:14087400:00011:00001",
  "USGS:14087400:00011:00002",
  "USGS:14087400:00011:00003",
  "USGS:14087520:00011:00001",
  "USGS:301124081395901:00011:00002",
  "USGS:301124081395901:00011:00006",
  "USGS:301124081395901:00011:00001",
  "USGS:301124081395901:00011:00005",
  "USGS:301124081395901:00011:00007",
  "USGS:301124081395901:00011:00009",
  "USGS:302309081333001:00011:00002",
  "USGS:302309081333001:00011:00006",
  "USGS:302309081333001:00011:00001",
  "USGS:302309081333001:00011:00005",
  "USGS:302309081333001:00011:00012",
  "USGS:302309081333001:00011:00014",
  "USGS:302309081333001:00011:00015",
  "USGS:302416081522601:00011:00002",
  "USGS:302847083145401:00011:00001",
  "USGS:303025085350501:00011:00002",
  "USGS:06442600:00011:00001",
  "USGS:06442996:00011:00003",
  "USGS:06445685:00011:00007",
  "USGS:06445685:00011:00002",
  "USGS:06445685:00011:00004",
  "USGS:06446000:00011:00002",
  "USGS:06446000:00011:00001",
  "USGS:06446500:00011:00004",
  "USGS:06446500:00011:00002",
  "USGS:06446500:00011:00005",
  "USGS:06446700:00011:00006",
  "USGS:06446700:00011:00002",
  "USGS:06446700:00011:00004",
  "USGS:06447230:00011:00005",
  "USGS:06447230:00011:00002",
  "USGS:06447230:00011:00004",
  "USGS:06447450:00011:00002",
  "USGS:06447450:00011:00004",
  "USGS:06447500:00011:00005",
  "USGS:06447500:00011:00001",
  "USGS:06447500:00011:00004",
  "USGS:06448000:00011:00001",
  "USGS:06448000:00011:00003",
  "USGS:02365500:00011:00002",
  "USGS:02365500:00011:00003",
  "USGS:02365769:00011:00002",
  "USGS:02365769:00011:00001",
  "USGS:02366000:00011:00001",
  "USGS:02366000:00011:00002",
  "USGS:02366500:00011:00002",
  "USGS:02366500:00011:00003",
  "USGS:02366650:00011:00002",
  "USGS:02366650:00011:00001",
  "USGS:02366996:00011:00002",
  "USGS:02366996:00011:00001",
  "USGS:02367310:00011:00002",
  "USGS:02367310:00011:00003",
  "USGS:02367900:00011:00002",
  "USGS:02367900:00011:00013",
  "USGS:02368000:00011:00002",
  "USGS:02368000:00011:00003",
  "USGS:02368500:00011:00001",
  "USGS:02368500:00011:00002",
  "USGS:02369000:00011:00003",
  "USGS:02369000:00011:00004",
  "USGS:02369600:00011:00018",
  "USGS:02369600:00011:00005",
  "USGS:02369600:00011:00004",
  "USGS:02370000:00011:00001",
  "USGS:02370000:00011:00002",
  "USGS:02370500:00011:00002",
  "USGS:02370500:00011:00003",
  "USGS:02375500:00011:00001",
  "USGS:02375500:00011:00005",
  "USGS:02376033:00011:00003",
  "USGS:02376033:00011:00001",
  "USGS:02376033:00011:00002",
  "USGS:02376100:00011:00003",
  "USGS:02376100:00011:00002",
  "USGS:02376115:00011:00002",
  "USGS:02376115:00011:00001",
  "USGS:02376293:00011:00002",
  "USGS:02376293:00011:00001",
  "USGS:250802081035500:00011:00014",
  "USGS:250802081035500:00011:00004",
  "USGS:250802081035500:00011:00005",
  "USGS:250802081035500:00011:00001",
  "USGS:250802081035500:00011:00002",
  "USGS:250802081035500:00011:00006",
  "USGS:250802081035500:00011:00008",
  "USGS:250802081035500:00011:00016",
  "USGS:250802081035500:00011:00030",
  "USGS:251003080435500:00011:00009",
  "USGS:251003080435500:00011:00012",
  "USGS:251003080435500:00011:00006",
  "USGS:251003080435500:00011:00033",
  "USGS:251003080435500:00011:00001",
  "USGS:251003080435500:00011:00008",
  "USGS:251003080435500:00011:00011",
  "USGS:251003080435500:00011:00024",
  "USGS:251003080435500:00011:00026",
  "USGS:251032080473400:00011:00003",
  "USGS:251032080473400:00011:00002",
  "USGS:251032080473400:00011:00001",
  "USGS:251115081075800:00011:00004",
  "USGS:251115081075800:00011:00005",
  "USGS:251115081075800:00011:00001",
  "USGS:251115081075800:00011:00002",
  "USGS:251115081075800:00011:00018",
  "USGS:251127080382100:00011:00009",
  "USGS:251127080382100:00011:00012",
  "USGS:251127080382100:00011:00026",
  "USGS:251127080382100:00011:00029",
  "USGS:251127080382100:00011:00030",
  "USGS:251127080382100:00011:00037",
  "USGS:251127080382100:00011:00001",
  "USGS:251127080382100:00011:00008",
  "USGS:251127080382100:00011:00011",
  "USGS:251127080382100:00011:00022",
  "USGS:251127080382100:00011:00024",
  "USGS:251209080350100:00011:00009",
  "USGS:251209080350100:00011:00012",
  "USGS:251209080350100:00011:00040",
  "USGS:251209080350100:00011:00001",
  "USGS:251209080350100:00011:00008",
  "USGS:251209080350100:00011:00011",
  "USGS:251209080350100:00011:00029",
  "USGS:251209080350100:00011:00031",
  "USGS:251241080385300:00011:00007",
  "USGS:251241080385300:00011:00008",
  "USGS:251241080385300:00011:00002",
  "USGS:251241080385300:00011:00003",
  "USGS:251241080385300:00011:00019",
  "USGS:251241080385300:00011:00001",
  "USGS:251241080385300:00011:00027",
  "USGS:251241080385300:00011:00028",
  "USGS:251241080385300:00011:00005",
  "USGS:251241080385300:00011:00006",
  "USGS:251253080320100:00011:00008",
  "USGS:251253080320100:00011:00009",
  "USGS:251253080320100:00011:00028",
  "USGS:251253080320100:00011:00037",
  "USGS:251253080320100:00011:00001",
  "USGS:251253080320100:00011:00005",
  "USGS:251253080320100:00011:00007",
  "USGS:251253080320100:00011:00024",
  "USGS:251253080320100:00011:00026",
  "USGS:251341080291200:00011:00008",
  "USGS:251341080291200:00011:00002",
  "USGS:251341080291200:00011:00003",
  "USGS:251341080291200:00011:00019",
  "USGS:251341080291200:00011:00001",
  "USGS:251341080291200:00011:00029",
  "USGS:251341080291200:00011:00006",
  "USGS:251355080312800:00011:00011",
  "USGS:251355080312800:00011:00041",
  "USGS:251355080312800:00011:00009",
  "USGS:251355080312800:00011:00012",
  "USGS:251355080312800:00011:00043",
  "USGS:251355080312800:00011:00022",
  "USGS:251355080312800:00011:00010",
  "USGS:251433080265000:00011:00008",
  "USGS:251433080265000:00011:00009",
  "USGS:251433080265000:00011:00039",
  "USGS:251433080265000:00011:00040",
  "USGS:251433080265000:00011:00032",
  "USGS:251433080265000:00011:00001",
  "USGS:251433080265000:00011:00005",
  "USGS:251433080265000:00011:00006",
  "USGS:251433080265000:00011:00023",
  "USGS:251433080265000:00011:00024",
  "USGS:251457080395802:00011:00001",
  "USGS:251457080395802:00011:00007",
  "USGS:251457080395802:00011:00016",
  "USGS:251457080395802:00011:00002",
  "USGS:251457080395802:00011:00005",
  "USGS:251457080395802:00011:00004",
  "USGS:251549080251200:00011:00015",
  "USGS:251549080251200:00011:00025",
  "USGS:251549080251200:00011:00043",
  "USGS:251549080251200:00011:00001",
  "USGS:251549080251200:00011:00024",
  "USGS:251549080251200:00011:00016",
  "USGS:251549080251200:00011:00017",
  "USGS:251549080251200:00011:00044",
  "USGS:251716080342100:00011:00001",
  "USGS:251716080342100:00011:00012",
  "USGS:251946080254800:00011:00001",
  "USGS:251946080254800:00011:00012",
  "USGS:252036080324300:00011:00001",
  "USGS:252230081021300:00011:00008",
  "USGS:252230081021300:00011:00002",
  "USGS:252230081021300:00011:00042",
  "USGS:252230081021300:00011:00001",
  "USGS:252230081021300:00011:00033",
  "USGS:252230081021300:00011:00006",
  "USGS:252230081021300:00011:00043",
  "USGS:252332080300501:00011:00001",
  "USGS:252502080253901:00011:00001",
  "USGS:252506080300601:00011:00010",
  "USGS:252551081050900:00011:00010",
  "USGS:252551081050900:00011:00013",
  "USGS:252551081050900:00011:00051",
  "USGS:252551081050900:00011:00017",
  "USGS:252551081050900:00011:00048",
  "USGS:252551081050900:00011:00053",
  "USGS:252551081050900:00011:00011",
  "USGS:252551081050900:00011:00012",
  "USGS:252551081050900:00011:00015",
  "USGS:252551081050900:00011:00035",
  "USGS:01133000:00011:00001",
  "USGS:01133000:00011:00002",
  "USGS:01134500:00011:00001",
  "USGS:01134500:00011:00003",
  "USGS:262724081260701:00011:00001",
  "USGS:262750080175001:00011:00001",
  "USGS:262750080175001:00011:00004",
  "USGS:263000080120001:00011:00001",
  "USGS:263000080120001:00011:00004",
  "USGS:263041081433102:00011:00001",
  "USGS:263041081433103:00011:00001",
  "USGS:263050080145001:00011:00001",
  "USGS:263050080145001:00011:00004",
  "USGS:263117082051001:00011:00001",
  "USGS:263117082051002:00011:00001",
  "USGS:263127081351602:00011:00001",
  "USGS:263180080205001:00011:00001",
  "USGS:263180080205001:00011:00004",
  "USGS:263251081452801:00011:00002",
  "USGS:263251081452802:00011:00002",
  "USGS:263251081452803:00011:00002",
  "USGS:263323081522401:00011:00001",
  "USGS:263335081394301:00011:00001",
  "USGS:263344081361703:00011:00001",
  "USGS:263440082022001:00011:00001",
  "USGS:263532081592201:00011:00001",
  "USGS:263537080211400:00011:00001",
  "USGS:263845081260701:00011:00001",
  "USGS:263845081260702:00011:00001",
  "USGS:263845081260703:00011:00001",
  "USGS:264053081572501:00011:00001",
  "USGS:264514080550700:00011:00021",
  "USGS:264514080550700:00011:00016",
  "USGS:264514080550700:00011:00017",
  "USGS:264755081460801:00011:00001",
  "USGS:264755081460802:00011:00001",
  "USGS:264941081321301:00011:00001",
  "USGS:265405080472100:00011:00016",
  "USGS:265405080472100:00011:00017",
  "USGS:265405080472100:00011:00018",
  "USGS:265405080472100:00011:00019",
  "USGS:265405080472100:00011:00020",
  "USGS:265405080472100:00011:00021",
  "USGS:265405080472100:00011:00022",
  "USGS:265405080472100:00011:00023",
  "USGS:265405080472100:00011:00024",
  "USGS:265405080472100:00011:00025",
  "USGS:265405080472100:00011:00013",
  "USGS:265405080472100:00011:00010",
  "USGS:265405080472100:00011:00012",
  "USGS:265405080472100:00011:00014",
  "USGS:265405080472100:00011:00009",
  "USGS:265405080472100:00011:00011",
  "USGS:265405080472100:00011:00008",
  "USGS:265405080472100:00011:00007",
  "USGS:265405080472100:00011:00006",
  "USGS:265405080472100:00011:00005",
  "USGS:265405080472100:00011:00004",
  "USGS:265501080364900:00011:00043",
  "USGS:265501080364900:00011:00016",
  "USGS:265501080364900:00011:00017",
  "USGS:265633080203001:00011:00001",
  "USGS:265651080045500:00011:00003",
  "USGS:14309000:00011:00003",
  "USGS:265651080045500:00011:00005",
  "USGS:265651080045500:00011:00001",
  "USGS:265651080045500:00011:00007",
  "USGS:265651080045500:00011:00008",
  "USGS:265651080045500:00011:00009",
  "USGS:265651080045500:00011:00010",
  "USGS:265812080053901:00011:00001",
  "USGS:265906080093500:00011:00011",
  "USGS:265906080093500:00011:00014",
  "USGS:265906080093500:00011:00001",
  "USGS:265906080093500:00011:00012",
  "USGS:265906080093500:00011:00015",
  "USGS:265906080093500:00011:00017",
  "USGS:265906080093500:00011:00018",
  "USGS:265929080091800:00011:00004",
  "USGS:265929080091800:00011:00001",
  "USGS:265929080091800:00011:00003",
  "USGS:265929080091800:00011:00005",
  "USGS:270124080280202:00011:00001",
  "USGS:270137082235301:00011:00002",
  "USGS:270157081203101:00011:00002",
  "USGS:270609080163401:00011:00001",
  "USGS:270835080105801:00011:00002",
  "USGS:270913080284901:00011:00001",
  "USGS:271538082002301:00011:00001",
  "USGS:271618080245801:00011:00001",
  "USGS:271619082240201:00011:00001",
  "USGS:271755080153001:00011:00002",
  "USGS:271755080153002:00011:00001",
  "USGS:271832082064801:00011:00001",
  "USGS:272012081482501:00011:00001",
  "USGS:05059310:00011:00002",
  "USGS:05059310:00011:00004",
  "USGS:05059480:00011:00002",
  "USGS:05059480:00011:00003",
  "USGS:05059500:00011:00004",
  "USGS:05059500:00011:00015",
  "USGS:05059600:00011:00002",
  "USGS:05059600:00011:00001",
  "USGS:05059700:00011:00001",
  "USGS:05059700:00011:00003",
  "USGS:05059715:00011:00007",
  "USGS:05059715:00011:00001",
  "USGS:05060000:00011:00001",
  "USGS:05060000:00011:00002",
  "USGS:05060100:00011:00002",
  "USGS:05060100:00011:00001",
  "USGS:05060100:00011:00008",
  "USGS:05060400:00011:00002",
  "USGS:05060500:00011:00001",
  "USGS:05060500:00011:00003",
  "USGS:05064500:00011:00006",
  "USGS:05064500:00011:00002",
  "USGS:05064500:00011:00005",
  "USGS:05064500:00011:00016",
  "USGS:05065500:00011:00001",
  "USGS:05065500:00011:00003",
  "USGS:05066500:00011:00001",
  "USGS:14161500:00011:00002",
  "USGS:14161500:00011:00003",
  "USGS:14162100:00011:00002",
  "USGS:14162200:00011:00001",
  "USGS:14162200:00011:00002",
  "USGS:14162200:00011:00003",
  "USGS:14162500:00011:00002",
  "USGS:14162500:00011:00003",
  "USGS:14162500:00011:00001",
  "USGS:14163150:00011:00002",
  "USGS:14163150:00011:00001",
  "USGS:14163900:00011:00002",
  "USGS:14163900:00011:00001",
  "USGS:14164550:00011:00001",
  "USGS:14164700:00011:00002",
  "USGS:14164700:00011:00001",
  "USGS:14164900:00011:00003",
  "USGS:14164900:00011:00002",
  "USGS:14165000:00011:00002",
  "USGS:14165000:00011:00003",
  "USGS:14165500:00011:00002",
  "USGS:14165500:00011:00003",
  "USGS:14166000:00011:00001",
  "USGS:14166000:00011:00002",
  "USGS:14166000:00011:00007",
  "USGS:14166500:00011:00001",
  "USGS:14166500:00011:00002",
  "USGS:14168000:00011:00002",
  "USGS:14169000:00011:00003",
  "USGS:14169000:00011:00001",
  "USGS:14169000:00011:00002",
  "USGS:14170000:00011:00001",
  "USGS:14170000:00011:00002",
  "USGS:14171000:00011:00001",
  "USGS:14171000:00011:00002",
  "USGS:14171600:00011:00002",
  "USGS:14171600:00011:00001",
  "USGS:14174000:00011:00003",
  "USGS:14174000:00011:00001",
  "USGS:14174000:00011:00002",
  "USGS:14178000:00011:00001",
  "USGS:14178000:00011:00002",
  "USGS:14178000:00011:00003",
  "USGS:14179000:00011:00001",
  "USGS:14179000:00011:00002",
  "USGS:14179000:00011:00003",
  "USGS:14180300:00011:00004",
  "USGS:14180300:00011:00002",
  "USGS:14180300:00011:00001",
  "USGS:14180500:00011:00003",
  "USGS:14180510:00011:00001",
  "USGS:14181400:00011:00001",
  "USGS:14181410:00011:00001",
  "USGS:14181500:00011:00001",
  "USGS:14181500:00011:00017",
  "USGS:14181500:00011:00015",
  "USGS:14181500:00011:00019",
  "USGS:14181500:00011:00002",
  "USGS:14181500:00011:00003",
  "USGS:14181500:00011:00005",
  "USGS:14181500:00011:00010",
  "USGS:14181500:00011:00008",
  "USGS:14181500:00011:00012",
  "USGS:14181500:00011:00006",
  "USGS:14181500:00011:00014",
  "USGS:14182500:00011:00001",
  "USGS:14182500:00011:00002",
  "USGS:14182500:00011:00003",
  "USGS:14182500:00011:00005",
  "USGS:14182500:00011:00011",
  "USGS:14182500:00011:00008",
  "USGS:14182500:00011:00006",
  "USGS:14183000:00011:00002",
  "USGS:14183000:00011:00003",
  "USGS:14183010:00011:00001",
  "USGS:14183010:00011:00002",
  "USGS:14183010:00011:00004",
  "USGS:14183010:00011:00005",
  "USGS:14184100:00011:00001",
  "USGS:14184100:00011:00002",
  "USGS:14184100:00011:00003",
  "USGS:14185000:00011:00002",
  "USGS:14185000:00011:00003",
  "USGS:14185000:00011:00004",
  "USGS:14185800:00011:00001",
  "USGS:14185800:00011:00003",
  "USGS:14185900:00011:00001",
  "USGS:14185900:00011:00002",
  "USGS:14185900:00011:00003",
  "USGS:14186100:00011:00002",
  "USGS:14186110:00011:00001",
  "USGS:14186200:00011:00001",
  "USGS:14186200:00011:00003",
  "USGS:14186600:00011:00002",
  "USGS:14186610:00011:00001",
  "USGS:06337000:00011:00025",
  "USGS:06337000:00011:00024",
  "USGS:06339100:00011:00001",
  "USGS:06339100:00011:00003",
  "USGS:06339500:00011:00002",
  "USGS:06339500:00011:00006",
  "USGS:06340000:00011:00001",
  "USGS:06340000:00011:00003",
  "USGS:06340500:00011:00002",
  "USGS:06340500:00011:00008",
  "USGS:06340700:00011:00004",
  "USGS:06341000:00011:00003",
  "USGS:06342020:00011:00003",
  "USGS:06342020:00011:00001",
  "USGS:06342260:00011:00001",
  "USGS:06342260:00011:00004",
  "USGS:06342450:00011:00001",
  "USGS:06342450:00011:00003",
  "USGS:06342500:00011:00001",
  "USGS:06342500:00011:00002",
  "USGS:06342500:00011:00007",
  "USGS:06342500:00011:00027",
  "USGS:06344600:00011:00001",
  "USGS:06344600:00011:00003",
  "USGS:06345500:00011:00001",
  "USGS:14190500:00011:00001",
  "USGS:14190500:00011:00002",
  "USGS:14191000:00011:00002",
  "USGS:14191000:00011:00003",
  "USGS:14192015:00011:00001",
  "USGS:14194150:00011:00002",
  "USGS:14194150:00011:00001",
  "USGS:14197900:00011:00003",
  "USGS:14197900:00011:00005",
  "USGS:14197900:00011:00002",
  "USGS:14197900:00011:00001",
  "USGS:14198400:00011:00002",
  "USGS:14198400:00011:00001",
  "USGS:14199704:00011:00002",
  "USGS:14199704:00011:00001",
  "USGS:14200000:00011:00002",
  "USGS:14200000:00011:00003",
  "USGS:14200100:00011:00002",
  "USGS:14200100:00011:00001",
  "USGS:14200300:00011:00004",
  "USGS:14200700:00011:00001",
  "USGS:14201300:00011:00001",
  "USGS:14201300:00011:00006",
  "USGS:14201300:00011:00002",
  "USGS:14201340:00011:00002",
  "USGS:14201340:00011:00001",
  "USGS:14201500:00011:00001",
  "USGS:14201500:00011:00002",
  "USGS:14202000:00011:00001",
  "USGS:14202000:00011:00002",
  "USGS:14309000:00011:00005",
  "USGS:14202630:00011:00001",
  "USGS:14202630:00011:00005",
  "USGS:14202980:00011:00003",
  "USGS:14202980:00011:00005",
  "USGS:14202980:00011:00006",
  "USGS:14202980:00011:00004",
  "USGS:14202980:00011:00007",
  "USGS:14203500:00011:00003",
  "USGS:14203500:00011:00001",
  "USGS:14205400:00011:00002",
  "USGS:14205400:00011:00001",
  "USGS:14206694:00011:00001",
  "USGS:14206694:00011:00004",
  "USGS:14206694:00011:00003",
  "USGS:14206694:00011:00002",
  "USGS:14206900:00011:00003",
  "USGS:14206900:00011:00002",
  "USGS:14206950:00011:00003",
  "USGS:14206950:00011:00002",
  "USGS:14206950:00011:00001",
  "USGS:14206950:00011:00004",
  "USGS:14206950:00011:00005",
  "USGS:14206950:00011:00006",
  "USGS:14206950:00011:00007",
  "USGS:14207200:00011:00001",
  "USGS:14207200:00011:00007",
  "USGS:14207200:00011:00009",
  "USGS:14207200:00011:00002",
  "USGS:14207200:00011:00003",
  "USGS:14207200:00011:00004",
  "USGS:14207500:00011:00003",
  "USGS:14207500:00011:00001",
  "USGS:14207740:00011:00002",
  "USGS:14207770:00011:00001",
  "USGS:14208700:00011:00001",
  "USGS:14208700:00011:00002",
  "USGS:14209000:00011:00007",
  "USGS:14209000:00011:00001",
  "USGS:14209000:00011:00002",
  "USGS:14209250:00011:00004",
  "USGS:14209250:00011:00001",
  "USGS:14209500:00011:00001",
  "USGS:14209500:00011:00003",
  "USGS:14209710:00011:00001",
  "USGS:14209710:00011:00002",
  "USGS:14209710:00011:00003",
  "USGS:14209710:00011:00004",
  "USGS:14209710:00011:00005",
  "USGS:14210000:00011:00004",
  "USGS:14210000:00011:00013",
  "USGS:14210000:00011:00001",
  "USGS:14210000:00011:00002",
  "USGS:14210000:00011:00007",
  "USGS:14210000:00011:00008",
  "USGS:14210000:00011:00009",
  "USGS:14210000:00011:00012",
  "USGS:14210000:00011:00010",
  "USGS:14211010:00011:00003",
  "USGS:14211010:00011:00002",
  "USGS:14211010:00011:00001",
  "USGS:14211010:00011:00004",
  "USGS:14211010:00011:00005",
  "USGS:14211010:00011:00006",
  "USGS:14211010:00011:00008",
  "USGS:14211010:00011:00007",
  "USGS:14211315:00011:00002",
  "USGS:14211315:00011:00001",
  "USGS:14211400:00011:00003",
  "USGS:14211400:00011:00002",
  "USGS:14211400:00011:00001",
  "USGS:14211499:00011:00003",
  "USGS:14211499:00011:00006",
  "USGS:14211499:00011:00002",
  "USGS:14211499:00011:00007",
  "USGS:14211499:00011:00001",
  "USGS:14211500:00011:00005",
  "USGS:14211500:00011:00001",
  "USGS:14211500:00011:00003",
  "USGS:14211550:00011:00003",
  "USGS:14211550:00011:00001",
  "USGS:14211550:00011:00002",
  "USGS:14211720:00011:00001",
  "USGS:14211720:00011:00005",
  "USGS:14211720:00011:00002",
  "USGS:14211720:00011:00003",
  "USGS:14211720:00011:00004",
  "USGS:14211720:00011:00036",
  "USGS:14211720:00011:00037",
  "USGS:14211720:00011:00039",
  "USGS:14211720:00011:00038",
  "USGS:14211720:00011:00041",
  "USGS:14211720:00011:00052",
  "USGS:14211720:00011:00055",
  "USGS:14211814:00011:00002",
  "USGS:14211814:00011:00001",
  "USGS:14211820:00011:00007",
  "USGS:14211820:00011:00003",
  "USGS:14211820:00011:00023",
  "USGS:14246900:00011:00023",
  "USGS:14246900:00011:00002",
  "USGS:14246900:00011:00003",
  "USGS:01142500:00011:00004",
  "USGS:01142500:00011:00001",
  "USGS:01142500:00011:00003",
  "USGS:01144000:00011:00001",
  "USGS:01144000:00011:00003",
  "USGS:01150900:00011:00005",
  "USGS:01150900:00011:00002",
  "USGS:01150900:00011:00003",
  "USGS:01151500:00011:00001",
  "USGS:01151500:00011:00004",
  "USGS:01153000:00011:00004",
  "USGS:01153000:00011:00003",
  "USGS:01153550:00011:00002",
  "USGS:01153550:00011:00006",
  "USGS:01154000:00011:00001",
  "USGS:01154000:00011:00002",
  "USGS:01155349:00011:00002",
  "USGS:01155349:00011:00001",
  "USGS:14301500:00011:00010",
  "USGS:14302020:00011:00003",
  "USGS:14302020:00011:00001",
  "USGS:14302480:00011:00004",
  "USGS:14302480:00011:00002",
  "USGS:14302480:00011:00001",
  "USGS:14302480:00011:00005",
  "USGS:14302480:00011:00009",
  "USGS:14302480:00011:00006",
  "USGS:14303200:00011:00001",
  "USGS:14303200:00011:00002",
  "USGS:14303200:00011:00004",
  "USGS:14303600:00011:00002",
  "USGS:14303600:00011:00003",
  "USGS:14305500:00011:00002",
  "USGS:14305500:00011:00003",
  "USGS:14306340:00011:00001",
  "USGS:14306340:00011:00006",
  "USGS:14306500:00011:00002",
  "USGS:14306500:00011:00006",
  "USGS:14307620:00011:00002",
  "USGS:14307620:00011:00006",
  "USGS:14308000:00011:00001",
  "USGS:14308000:00011:00002",
  "USGS:14308500:00011:00001",
  "USGS:14308500:00011:00002",
  "USGS:14308990:00011:00001",
  "USGS:14308990:00011:00004",
  "USGS:14308995:00011:00001",
  "USGS:14309000:00011:00002",
  "USGS:14309500:00011:00001",
  "USGS:14309500:00011:00003",
  "USGS:14310000:00011:00001",
  "USGS:14310000:00011:00002",
  "USGS:14312000:00011:00001",
  "USGS:14312000:00011:00003",
  "USGS:14312450:00011:00001",
  "USGS:14312500:00011:00001",
  "USGS:14312500:00011:00002",
  "USGS:14313000:00011:00001",
  "USGS:14313200:00011:00002",
  "USGS:14313200:00011:00001",
  "USGS:14313500:00011:00001",
  "USGS:14313500:00011:00002",
  "USGS:14313700:00011:00002",
  "USGS:14313700:00011:00001",
  "USGS:14314500:00011:00001",
  "USGS:14314500:00011:00002",
  "USGS:14314700:00011:00002",
  "USGS:14314700:00011:00001",
  "USGS:14315500:00011:00001",
  "USGS:14315500:00011:00002",
  "USGS:14315700:00011:00002",
  "USGS:14315700:00011:00001",
  "USGS:14315950:00011:00002",
  "USGS:14315950:00011:00001",
  "USGS:14316455:00011:00002",
  "USGS:14316455:00011:00001",
  "USGS:14316460:00011:00003",
  "USGS:14316460:00011:00001",
  "USGS:14316460:00011:00004",
  "USGS:14316460:00011:00002",
  "USGS:14316460:00011:00005",
  "USGS:14316495:00011:00004",
  "USGS:14316495:00011:00002",
  "USGS:14316495:00011:00001",
  "USGS:14316500:00011:00005",
  "USGS:14316500:00011:00001",
  "USGS:14316500:00011:00002",
  "USGS:14316500:00011:00007",
  "USGS:14316700:00011:00001",
  "USGS:14316700:00011:00002",
  "USGS:14317450:00011:00003",
  "USGS:14317450:00011:00001",
  "USGS:14317450:00011:00004",
  "USGS:14317450:00011:00002",
  "USGS:14317450:00011:00005",
  "USGS:14318000:00011:00003",
  "USGS:14318000:00011:00001",
  "USGS:14318000:00011:00002",
  "USGS:14319500:00011:00002",
  "USGS:14319500:00011:00003",
  "USGS:14320934:00011:00002",
  "USGS:14320934:00011:00003",
  "USGS:14320934:00011:00001",
  "USGS:14321000:00011:00002",
  "USGS:14321000:00011:00003",
  "USGS:14325000:00011:00001",
  "USGS:14325000:00011:00002",
  "USGS:14326510:00011:00001",
  "USGS:14327000:00011:00002",
  "USGS:14327055:00011:00001",
  "USGS:14330000:00011:00001",
  "USGS:14330000:00011:00002",
  "USGS:14330000:00011:00003",
  "USGS:14332000:00011:00001",
  "USGS:14332000:00011:00002",
  "USGS:14335040:00011:00001",
  "USGS:14335072:00011:00003",
  "USGS:14335072:00011:00001",
  "USGS:14335072:00011:00002",
  "USGS:14337500:00011:00003",
  "USGS:14337500:00011:00004",
  "USGS:14337600:00011:00001",
  "USGS:14337600:00011:00002",
  "USGS:14337600:00011:00003",
  "USGS:01613900:00011:00001",
  "USGS:01613900:00011:00005",
  "USGS:01615000:00011:00001",
  "USGS:01615000:00011:00002",
  "USGS:01616100:00011:00004",
  "USGS:01616100:00011:00002",
  "USGS:01616100:00011:00001",
  "USGS:01616100:00011:00005",
  "USGS:01620500:00011:00001",
  "USGS:01620500:00011:00005",
  "USGS:01621050:00011:00002",
  "USGS:01621050:00011:00003",
  "USGS:01622000:00011:00001",
  "USGS:06409000:00011:00002",
  "USGS:06409000:00011:00008",
  "USGS:06410000:00011:00001",
  "USGS:06410000:00011:00006",
  "USGS:06410500:00011:00005",
  "USGS:06410500:00011:00001",
  "USGS:06410500:00011:00003",
  "USGS:06411500:00011:00002",
  "USGS:06411500:00011:00007",
  "USGS:06412500:00011:00006",
  "USGS:06412500:00011:00002",
  "USGS:06412500:00011:00005",
  "USGS:06412810:00011:00002",
  "USGS:06412810:00011:00006",
  "USGS:06414000:00011:00005",
  "USGS:06414000:00011:00001",
  "USGS:06414000:00011:00003",
  "USGS:06418900:00011:00010",
  "USGS:06418900:00011:00001",
  "USGS:06418900:00011:00007",
  "USGS:06421500:00011:00005",
  "USGS:06421500:00011:00002",
  "USGS:06421500:00011:00003",
  "USGS:06422500:00011:00008",
  "USGS:06422500:00011:00002",
  "USGS:06422500:00011:00006",
  "USGS:06423500:00011:00001",
  "USGS:06423500:00011:00006",
  "USGS:06423500:00011:00003",
  "USGS:06424000:00011:00009",
  "USGS:06424000:00011:00002",
  "USGS:06424000:00011:00007",
  "USGS:06425100:00011:00006",
  "USGS:06425100:00011:00001",
  "USGS:06425100:00011:00004",
  "USGS:06425500:00011:00006",
  "USGS:06425500:00011:00001",
  "USGS:06425500:00011:00004",
  "USGS:06428500:00011:00007",
  "USGS:06428500:00011:00002",
  "USGS:06428500:00011:00005",
  "USGS:06429997:00011:00001",
  "USGS:06429997:00011:00004",
  "USGS:06430500:00011:00008",
  "USGS:06430500:00011:00001",
  "USGS:06430500:00011:00006",
  "USGS:06430532:00011:00002",
  "USGS:06430532:00011:00003",
  "USGS:06430770:00011:00002",
  "USGS:06430770:00011:00003",
  "USGS:06430800:00011:00008",
  "USGS:06430800:00011:00002",
  "USGS:06430800:00011:00007",
  "USGS:06430850:00011:00002",
  "USGS:06430850:00011:00004",
  "USGS:06431500:00011:00006",
  "USGS:06431500:00011:00001",
  "USGS:06431500:00011:00004",
  "USGS:06433000:00011:00009",
  "USGS:06433000:00011:00001",
  "USGS:06433000:00011:00007",
  "USGS:06434505:00011:00005",
  "USGS:06434505:00011:00002",
  "USGS:06434505:00011:00007",
  "USGS:06436000:00011:00007",
  "USGS:06436000:00011:00001",
  "USGS:06436000:00011:00004",
  "USGS:06436165:00011:00004",
  "USGS:06436165:00011:00002",
  "USGS:06436165:00011:00001",
  "USGS:06436180:00011:00008",
  "USGS:06436180:00011:00001",
  "USGS:06436180:00011:00006",
  "USGS:06436190:00011:00007",
  "USGS:06436190:00011:00001",
  "USGS:06436190:00011:00004",
  "USGS:06436198:00011:00001",
  "USGS:06436198:00011:00004",
  "USGS:06437000:00011:00007",
  "USGS:06437000:00011:00002",
  "USGS:06437000:00011:00005",
  "USGS:06437020:00011:00002",
  "USGS:06437020:00011:00004",
  "USGS:06438000:00011:00007",
  "USGS:06438000:00011:00002",
  "USGS:06438000:00011:00005",
  "USGS:06438500:00011:00016",
  "USGS:06438500:00011:00014",
  "USGS:06438500:00011:00001",
  "USGS:06438500:00011:00015",
  "USGS:06440000:00011:00016",
  "USGS:06440000:00011:00013",
  "USGS:06440200:00011:00010",
  "USGS:06440200:00011:00002",
  "USGS:06440200:00011:00009",
  "USGS:06441500:00011:00004",
  "USGS:06441500:00011:00007",
  "USGS:06441500:00011:00002",
  "USGS:06441590:00011:00002",
  "USGS:06441592:00011:00001",
  "USGS:06441595:00011:00002",
  "USGS:06442130:00011:00004",
  "USGS:350624081023345:00011:00004",
  "USGS:02136000:00011:00018",
  "USGS:02136000:00011:00001",
  "USGS:02136000:00011:00002",
  "USGS:02136361:00011:00011",
  "USGS:02136361:00011:00001",
  "USGS:021457492:00011:00003",
  "USGS:021457492:00011:00001",
  "USGS:021459367:00011:00003",
  "USGS:021459367:00011:00001",
  "USGS:02146000:00011:00009",
  "USGS:02146000:00011:00008",
  "USGS:02146110:00011:00003",
  "USGS:02146110:00011:00001",
  "USGS:0214676115:00011:00002",
  "USGS:0214676115:00011:00001",
  "USGS:02146800:00011:00003",
  "USGS:02146800:00011:00002",
  "USGS:02147020:00011:00015",
  "USGS:06400875:00011:00005",
  "USGS:06401500:00011:00006",
  "USGS:06401500:00011:00005",
  "USGS:06401500:00011:00002",
  "USGS:06402000:00011:00005",
  "USGS:06402000:00011:00004",
  "USGS:06402000:00011:00002",
  "USGS:06402430:00011:00002",
  "USGS:06402430:00011:00003",
  "USGS:06402500:00011:00010",
  "USGS:06402500:00011:00001",
  "USGS:06402500:00011:00009",
  "USGS:06402600:00011:00002",
  "USGS:06402600:00011:00001",
  "USGS:06403300:00011:00001",
  "USGS:06403300:00011:00003",
  "USGS:09180000:00011:00001",
  "USGS:09180000:00011:00002",
  "USGS:09180000:00011:00003",
  "USGS:09180000:00011:00004",
  "USGS:09180000:00011:00013",
  "USGS:09180500:00011:00001",
  "USGS:09180500:00011:00003",
  "USGS:09180500:00011:00004",
  "USGS:09180500:00011:00005",
  "USGS:09182400:00011:00002",
  "USGS:09182400:00011:00001",
  "USGS:14338000:00011:00005",
  "USGS:14338000:00011:00001",
  "USGS:14338000:00011:00002",
  "USGS:14338000:00011:00007",
  "USGS:14339000:00011:00005",
  "USGS:14339000:00011:00006",
  "USGS:14339000:00011:00001",
  "USGS:14353000:00011:00001",
  "USGS:14353000:00011:00002",
  "USGS:14353500:00011:00001",
  "USGS:14353500:00011:00002",
  "USGS:14354200:00011:00002",
  "USGS:14354200:00011:00001",
  "USGS:14354200:00011:00004",
  "USGS:14354200:00011:00003",
  "USGS:14357500:00011:00001",
  "USGS:14357500:00011:00002",
  "USGS:14359000:00011:00017",
  "USGS:14359000:00011:00006",
  "USGS:14359000:00011:00001",
  "USGS:14361500:00011:00005",
  "USGS:14361500:00011:00006",
  "USGS:14361500:00011:00007",
  "USGS:14361500:00011:00018",
  "USGS:14361900:00011:00003",
  "USGS:14362000:00011:00003",
  "USGS:14362000:00011:00006",
  "USGS:14362000:00011:00002",
  "USGS:14362250:00011:00001",
  "USGS:14362250:00011:00002",
  "USGS:14366000:00011:00015",
  "USGS:14366000:00011:00005",
  "USGS:14366000:00011:00002",
  "USGS:14369500:00011:00003",
  "USGS:14369500:00011:00001",
  "USGS:14369500:00011:00002",
  "USGS:14372300:00011:00001",
  "USGS:14372300:00011:00002",
  "USGS:14372300:00011:00004",
  "USGS:14375100:00011:00001",
  "USGS:14375100:00011:00002",
  "USGS:14377100:00011:00001",
  "USGS:14377100:00011:00002",
  "USGS:14400000:00011:00001",
  "USGS:14400000:00011:00004",
  "USGS:420451121510000:00011:00001",
  "USGS:420451121510000:00011:00004",
  "USGS:420451121510000:00011:00005",
  "USGS:420451121510000:00011:00002",
  "USGS:420451121510000:00011:00003",
  "USGS:420741121554001:00011:00001",
  "USGS:420741121554001:00011:00004",
  "USGS:420741121554001:00011:00005",
  "USGS:420741121554001:00011:00002",
  "USGS:420741121554001:00011:00003",
  "USGS:420853121505500:00011:00001",
  "USGS:420853121505500:00011:00004",
  "USGS:420853121505500:00011:00005",
  "USGS:420853121505500:00011:00002",
  "USGS:420853121505500:00011:00003",
  "USGS:420853121505501:00011:00001",
  "USGS:420853121505501:00011:00004",
  "USGS:420853121505501:00011:00005",
  "USGS:420853121505501:00011:00002",
  "USGS:420853121505501:00011:00003",
  "USGS:421015121471800:00011:00001",
  "USGS:421015121471800:00011:00004",
  "USGS:421015121471800:00011:00005",
  "USGS:421015121471800:00011:00002",
  "USGS:421015121471800:00011:00003",
  "USGS:421401121480900:00011:00001",
  "USGS:421401121480900:00011:00004",
  "USGS:421401121480900:00011:00005",
  "USGS:421401121480900:00011:00002",
  "USGS:421401121480900:00011:00003",
  "USGS:434400121275801:00011:00001",
  "USGS:442242121405501:00011:00001",
  "USGS:452033122195901:00011:00001",
  "USGS:452359122454500:00011:00005",
  "USGS:452359122454500:00011:00001",
  "USGS:452912122312801:00011:00001",
  "USGS:452912122312801:00011:00003",
  "USGS:453004122510301:00011:00001",
  "USGS:453004122510301:00011:00003",
  "USGS:453004122510301:00011:00004",
  "USGS:453004122510301:00011:00002",
  "USGS:453004122510301:00011:00006",
  "USGS:453030122560101:00011:00001",
  "USGS:453030122560101:00011:00003",
  "USGS:453030122560101:00011:00004",
  "USGS:453030122560101:00011:00002",
  "USGS:453030122560101:00011:00006",
  "USGS:453040123065201:00011:00001",
  "USGS:453040123065201:00011:00003",
  "USGS:453040123065201:00011:00004",
  "USGS:453040123065201:00011:00002",
  "USGS:453040123065201:00011:00006",
  "USGS:453630122021400:00011:00014",
  "USGS:453630122021400:00011:00015",
  "USGS:453630122021400:00011:00016",
  "USGS:453630122021400:00011:00005",
  "USGS:453630122021400:00011:00018",
  "USGS:455009119142301:00011:00001",
  "USGS:455009119142301:00011:00002",
  "USGS:455009119142301:00011:00004",
  "USGS:455009119142301:00011:00003",
  "USGS:455415119314601:00011:00001",
  "USGS:455415119314601:00011:00002",
  "USGS:455415119314601:00011:00004",
  "USGS:455415119314601:00011:00003",
  "USGS:02163500:00011:00016",
  "USGS:02163500:00011:00015",
  "USGS:02164000:00011:00017",
  "USGS:02164000:00011:00001",
  "USGS:02164000:00011:00002",
  "USGS:02164110:00011:00015",
  "USGS:02164110:00011:00005",
  "USGS:021650905:00011:00003",
  "USGS:021650905:00011:00001",
  "USGS:01135150:00011:00002",
  "USGS:01135150:00011:00003",
  "USGS:01135300:00011:00002",
  "USGS:01135300:00011:00003",
  "USGS:01135500:00011:00001",
  "USGS:01135500:00011:00003",
  "USGS:01138500:00011:00002",
  "USGS:01138500:00011:00005",
  "USGS:01139000:00011:00001",
  "USGS:01139000:00011:00004",
  "USGS:01139800:00011:00004",
  "USGS:01139800:00011:00001",
  "USGS:01139800:00011:00003",
  "USGS:01141500:00011:00006",
  "USGS:01141500:00011:00005",
  "USGS:06480000:00011:00019",
  "USGS:06480000:00011:00010",
  "USGS:06480000:00011:00001",
  "USGS:06480000:00011:00009",
  "USGS:06481000:00011:00006",
  "USGS:06481000:00011:00002",
  "USGS:06481000:00011:00004",
  "USGS:06481400:00011:00004",
  "USGS:06481400:00011:00001",
  "USGS:06481480:00011:00004",
  "USGS:06481480:00011:00001",
  "USGS:06481480:00011:00003",
  "USGS:06481493:00011:00001",
  "USGS:06481497:00011:00001",
  "USGS:06481500:00011:00005",
  "USGS:06481500:00011:00001",
  "USGS:06481500:00011:00003",
  "USGS:06482000:00011:00003",
  "USGS:06482000:00011:00001",
  "USGS:06482000:00011:00002",
  "USGS:06482010:00011:00001",
  "USGS:06482020:00011:00001",
  "USGS:06482020:00011:00007",
  "USGS:06482020:00011:00003",
  "USGS:06482610:00011:00005",
  "USGS:06482610:00011:00001",
  "USGS:06482610:00011:00003",
  "USGS:430027102311801:00011:00001",
  "USGS:430027102311806:00011:00006",
  "USGS:430027102311806:00011:00001",
  "USGS:430314100372001:00011:00004",
  "USGS:430314100372001:00011:00003",
  "USGS:430337100243201:00011:00004",
  "USGS:430337100243201:00011:00001",
  "USGS:430415100451501:00011:00004",
  "USGS:430415100451501:00011:00003",
  "USGS:430726101033501:00011:00004",
  "USGS:430726101033501:00011:00001",
  "USGS:431158100461002:00011:00003",
  "USGS:431158100461002:00011:00001",
  "USGS:431428100192701:00011:00004",
  "USGS:431428100192701:00011:00001",
  "USGS:433047096391700:00011:00001",
  "USGS:433141096572100:00011:00001",
  "USGS:433326096405200:00011:00001",
  "USGS:433600096442400:00011:00001",
  "USGS:433726096444501:00011:00001",
  "USGS:433752096432701:00011:00001",
  "USGS:434329096521201:00011:00001",
  "USGS:434330096434801:00011:00002",
  "USGS:434913097041800:00011:00001",
  "USGS:440326103180702:00011:00002",
  "USGS:440544103180001:00011:00001",
  "USGS:440544103180002:00011:00001",
  "USGS:441759103261202:00011:00002",
  "USGS:441759103261202:00011:00001",
  "USGS:441759103261203:00011:00003",
  "USGS:445959096582600:00011:00001",
  "USGS:450628097060800:00011:00001",
  "USGS:451605097071701:00011:00002",
  "USGS:451605097071701:00011:00001",
  "USGS:452115097110601:00011:00003",
  "USGS:452304097083901:00011:00001",
  "USGS:453358098260101:00011:00001",
  "USGS:453515097083801:00011:00003",
  "USGS:453819096572501:00011:00004",
  "USGS:453819096572501:00011:00001",
  "USGS:021720677:00011:00002",
  "USGS:021720677:00011:00001",
  "USGS:021720677:00011:00003",
  "USGS:021720677:00011:00004",
  "USGS:02147020:00011:00005",
  "USGS:021473415:00011:00003",
  "USGS:021473415:00011:00001",
  "USGS:021473426:00011:00005",
  "USGS:021473426:00011:00001",
  "USGS:021473428:00011:00005",
  "USGS:021473428:00011:00001",
  "USGS:02147500:00011:00001",
  "USGS:02147500:00011:00002",
  "USGS:02148000:00011:00016",
  "USGS:02148000:00011:00001",
  "USGS:02148000:00011:00002",
  "USGS:02153051:00011:00001",
  "USGS:02153200:00011:00011",
  "USGS:02153200:00011:00001",
  "USGS:02153500:00011:00004",
  "USGS:02153500:00011:00001",
  "USGS:02153500:00011:00002",
  "USGS:02153525:00011:00003",
  "USGS:02153525:00011:00002",
  "USGS:02153550:00011:00003",
  "USGS:02153551:00011:00003",
  "USGS:02153551:00011:00001",
  "USGS:02153590:00011:00002",
  "USGS:02153590:00011:00001",
  "USGS:02153700:00011:00002",
  "USGS:02153700:00011:00001",
  "USGS:02154500:00011:00014",
  "USGS:02154500:00011:00004",
  "USGS:02154790:00011:00014",
  "USGS:02154790:00011:00004",
  "USGS:02154950:00011:00001",
  "USGS:02155500:00011:00015",
  "USGS:02155500:00011:00005",
  "USGS:02155500:00011:00004",
  "USGS:021556524:00011:00003",
  "USGS:021556525:00011:00013",
  "USGS:021556525:00011:00001",
  "USGS:02156300:00011:00006",
  "USGS:02156300:00011:00003",
  "USGS:02156449:00011:00003",
  "USGS:021564493:00011:00002",
  "USGS:021564493:00011:00001",
  "USGS:02156500:00011:00003",
  "USGS:02156500:00011:00005",
  "USGS:02156500:00011:00006",
  "USGS:02156500:00011:00001",
  "USGS:02156500:00011:00002",
  "USGS:02156500:00011:00004",
  "USGS:02157470:00011:00002",
  "USGS:02157470:00011:00001",
  "USGS:02157510:00011:00002",
  "USGS:02157510:00011:00001",
  "USGS:02158408:00011:00002",
  "USGS:02158408:00011:00001",
  "USGS:02160105:00011:00003",
  "USGS:02160105:00011:00005",
  "USGS:02160105:00011:00006",
  "USGS:02160105:00011:00001",
  "USGS:02160105:00011:00002",
  "USGS:02160105:00011:00004",
  "USGS:02160325:00011:00003",
  "USGS:02160325:00011:00001",
  "USGS:02160326:00011:00011",
  "USGS:02160326:00011:00001",
  "USGS:02160381:00011:00013",
  "USGS:02160381:00011:00011",
  "USGS:02160381:00011:00001",
  "USGS:02160390:00011:00011",
  "USGS:02160390:00011:00001",
  "USGS:02160700:00011:00003",
  "USGS:02160700:00011:00005",
  "USGS:02160700:00011:00006",
  "USGS:02160700:00011:00001",
  "USGS:02160700:00011:00002",
  "USGS:02160700:00011:00004",
  "USGS:02160990:00011:00003",
  "USGS:02160991:00011:00003",
  "USGS:02160991:00011:00032",
  "USGS:02160991:00011:00001",
  "USGS:02160991:00011:00002",
  "USGS:02160991:00011:00004",
  "USGS:02161000:00011:00001",
  "USGS:02161000:00011:00002",
  "USGS:02162035:00011:00003",
  "USGS:02162035:00011:00002",
  "USGS:02162035:00011:00012",
  "USGS:02162035:00011:00001",
  "USGS:02162035:00011:00004",
  "USGS:02162035:00011:00005",
  "USGS:02162035:00011:00006",
  "USGS:02162093:00011:00001",
  "USGS:02162093:00011:00002",
  "USGS:02162290:00011:00002",
  "USGS:02162290:00011:00001",
  "USGS:02162350:00011:00004",
  "USGS:02162500:00011:00004",
  "USGS:02162500:00011:00003",
  "USGS:02163001:00011:00001",
  "USGS:02163001:00011:00012",
  "USGS:02163001:00011:00002",
  "USGS:01442500:00011:00004",
  "USGS:01442500:00011:00003",
  "USGS:01446775:00011:00002",
  "USGS:01446775:00011:00001",
  "USGS:01447500:00011:00003",
  "USGS:01447500:00011:00004",
  "USGS:01447500:00011:00001",
  "USGS:01447500:00011:00002",
  "USGS:01447680:00011:00004",
  "USGS:01447680:00011:00003",
  "USGS:01447720:00011:00003",
  "USGS:01447720:00011:00004",
  "USGS:01447720:00011:00001",
  "USGS:01447720:00011:00002",
  "USGS:01447780:00011:00002",
  "USGS:01447780:00011:00001",
  "USGS:01447800:00011:00003",
  "USGS:01447800:00011:00001",
  "USGS:01447800:00011:00002",
  "USGS:01449000:00011:00003",
  "USGS:06449000:00011:00001",
  "USGS:06449000:00011:00004",
  "USGS:06449100:00011:00001",
  "USGS:06449100:00011:00006",
  "USGS:06449500:00011:00001",
  "USGS:06449500:00011:00009",
  "USGS:06450500:00011:00006",
  "USGS:06450500:00011:00002",
  "USGS:06450500:00011:00003",
  "USGS:06452000:00011:00001",
  "USGS:06452000:00011:00006",
  "USGS:06452000:00011:00018",
  "USGS:06452320:00011:00006",
  "USGS:06452320:00011:00002",
  "USGS:06452320:00011:00004",
  "USGS:06453020:00011:00002",
  "USGS:06464100:00011:00009",
  "USGS:06464100:00011:00001",
  "USGS:06464100:00011:00006",
  "USGS:06464500:00011:00009",
  "USGS:06464500:00011:00001",
  "USGS:06464500:00011:00007",
  "USGS:06466700:00011:00013",
  "USGS:06466700:00011:00001",
  "USGS:06467500:00011:00021",
  "USGS:06467500:00011:00001",
  "USGS:06467500:00011:00003",
  "USGS:06470878:00011:00005",
  "USGS:06470878:00011:00002",
  "USGS:06470878:00011:00006",
  "USGS:06471000:00011:00002",
  "USGS:06471000:00011:00007",
  "USGS:06471065:00011:00004",
  "USGS:06471065:00011:00001",
  "USGS:06471500:00011:00011",
  "USGS:06471500:00011:00003",
  "USGS:06471500:00011:00008",
  "USGS:06471510:00011:00004",
  "USGS:06471510:00011:00001",
  "USGS:06471770:00011:00001",
  "USGS:06471800:00011:00004",
  "USGS:06471800:00011:00002",
  "USGS:06471800:00011:00001",
  "USGS:06472000:00011:00005",
  "USGS:06472000:00011:00001",
  "USGS:06472000:00011:00003",
  "USGS:06473000:00011:00019",
  "USGS:06473000:00011:00002",
  "USGS:06473000:00011:00008",
  "USGS:06475000:00011:00015",
  "USGS:06475000:00011:00002",
  "USGS:06475000:00011:00004",
  "USGS:06476000:00011:00023",
  "USGS:06476000:00011:00002",
  "USGS:06476000:00011:00007",
  "USGS:06477000:00011:00005",
  "USGS:06477000:00011:00001",
  "USGS:06477000:00011:00004",
  "USGS:06477500:00011:00006",
  "USGS:06477500:00011:00001",
  "USGS:06477500:00011:00004",
  "USGS:06478000:00011:00002",
  "USGS:06478000:00011:00001",
  "USGS:06478500:00011:00001",
  "USGS:06478500:00011:00006",
  "USGS:06478500:00011:00003",
  "USGS:06478513:00011:00003",
  "USGS:06478513:00011:00006",
  "USGS:06478600:00011:00002",
  "USGS:06478600:00011:00003",
  "USGS:06478690:00011:00009",
  "USGS:06478690:00011:00001",
  "USGS:06478690:00011:00007",
  "USGS:06479010:00011:00018",
  "USGS:06479010:00011:00001",
  "USGS:06479010:00011:00005",
  "USGS:06479010:00011:00003",
  "USGS:06479215:00011:00015",
  "USGS:06479215:00011:00001",
  "USGS:06479215:00011:00003",
  "USGS:06479438:00011:00018",
  "USGS:06479438:00011:00001",
  "USGS:06479438:00011:00003",
  "USGS:06479449:00011:00001",
  "USGS:06479490:00011:00006",
  "USGS:06479490:00011:00003",
  "USGS:06479498:00011:00004",
  "USGS:06479498:00011:00001",
  "USGS:06479500:00011:00003",
  "USGS:06479500:00011:00001",
  "USGS:06479500:00011:00002",
  "USGS:06479512:00011:00001",
  "USGS:06479515:00011:00003",
  "USGS:06479525:00011:00016",
  "USGS:06479525:00011:00001",
  "USGS:06479525:00011:00003",
  "USGS:06479770:00011:00005",
  "USGS:06479770:00011:00002",
  "USGS:06479770:00011:00004",
  "USGS:01519995:00011:00013",
  "USGS:01519995:00011:00002",
  "USGS:01519995:00011:00001",
  "USGS:01520000:00011:00003",
  "USGS:01520000:00011:00001",
  "USGS:01520000:00011:00002",
  "USGS:01531250:00011:00001",
  "USGS:01531250:00011:00002",
  "USGS:01531325:00011:00002",
  "USGS:01531325:00011:00001",
  "USGS:01531500:00011:00001",
  "USGS:01531500:00011:00002",
  "USGS:01531908:00011:00002",
  "USGS:01531908:00011:00001",
  "USGS:01532000:00011:00004",
  "USGS:01532000:00011:00003",
  "USGS:01533400:00011:00004",
  "USGS:01533400:00011:00003",
  "USGS:01534000:00011:00007",
  "USGS:01534000:00011:00006",
  "USGS:01534000:00011:00005",
  "USGS:01534180:00011:00013",
  "USGS:01534180:00011:00002",
  "USGS:06345500:00011:00005",
  "USGS:06345780:00011:00002",
  "USGS:06345780:00011:00004",
  "USGS:06347000:00011:00001",
  "USGS:06347000:00011:00003",
  "USGS:06347500:00011:00001",
  "USGS:06347500:00011:00003",
  "USGS:06348300:00011:00004",
  "USGS:06348300:00011:00001",
  "USGS:06348500:00011:00001",
  "USGS:06348500:00011:00002",
  "USGS:06349000:00011:00002",
  "USGS:06349000:00011:00008",
  "USGS:06349070:00011:00001",
  "USGS:06349070:00011:00002",
  "USGS:06349070:00011:00013",
  "USGS:06349070:00011:00014",
  "USGS:06349500:00011:00001",
  "USGS:06349500:00011:00003",
  "USGS:06349600:00011:00002",
  "USGS:06349600:00011:00001",
  "USGS:06349700:00011:00004",
  "USGS:06349700:00011:00001",
  "USGS:06350000:00011:00002",
  "USGS:06350000:00011:00007",
  "USGS:06351200:00011:00015",
  "USGS:06351200:00011:00014",
  "USGS:06352000:00011:00001",
  "USGS:06352000:00011:00003",
  "USGS:06353000:00011:00001",
  "USGS:06353000:00011:00003",
  "USGS:06354000:00011:00002",
  "USGS:06354000:00011:00007",
  "USGS:06354480:00011:00004",
  "USGS:06354480:00011:00001",
  "USGS:06354490:00011:00001",
  "USGS:06354580:00011:00002",
  "USGS:06354580:00011:00003",
  "USGS:06468170:00011:00001",
  "USGS:06468170:00011:00007",
  "USGS:06468250:00011:00001",
  "USGS:06468250:00011:00006",
  "USGS:06469400:00011:00001",
  "USGS:06469400:00011:00003",
  "USGS:06470000:00011:00001",
  "USGS:06470000:00011:00007",
  "USGS:06470500:00011:00002",
  "USGS:06470500:00011:00005",
  "USGS:06470800:00011:00001",
  "USGS:06470800:00011:00003",
  "USGS:06471200:00011:00006",
  "USGS:06471200:00011:00001",
  "USGS:06471200:00011:00004",
  "USGS:460120097591803:00011:00001",
  "USGS:461838097553402:00011:00001",
  "USGS:462400097552502:00011:00001",
  "USGS:462425096441202:00011:00001",
  "USGS:462633097163402:00011:00001",
  "USGS:463417099271002:00011:00001",
  "USGS:463422097115602:00011:00001",
  "USGS:464114097260900:00011:00002",
  "USGS:464114097260900:00011:00001",
  "USGS:464114097260900:00011:00006",
  "USGS:464114097260900:00011:00007",
  "USGS:464114097260900:00011:00008",
  "USGS:464114097260900:00011:00009",
  "USGS:464114097260900:00011:00005",
  "USGS:464115097254700:00011:00002",
  "USGS:464115097254700:00011:00001",
  "USGS:464115097255000:00011:00004",
  "USGS:464115097255000:00011:00008",
  "USGS:464115097255000:00011:00009",
  "USGS:464115097255000:00011:00013",
  "USGS:464115097255000:00011:00005",
  "USGS:464115097255000:00011:00002",
  "USGS:464115097255000:00011:00001",
  "USGS:464540100222101:00011:00001",
  "USGS:464703100464600:00011:00001",
  "USGS:01470960:00011:00003",
  "USGS:01470960:00011:00001",
  "USGS:01470960:00011:00002",
  "USGS:01471000:00011:00001",
  "USGS:01471000:00011:00002",
  "USGS:01471510:00011:00003",
  "USGS:01471510:00011:00001",
  "USGS:01471510:00011:00002",
  "USGS:01471875:00011:00004",
  "USGS:01471875:00011:00003",
  "USGS:05066500:00011:00003",
  "USGS:05070000:00011:00002",
  "USGS:05070000:00011:00001",
  "USGS:05082500:00011:00024",
  "USGS:05082500:00011:00002",
  "USGS:05082500:00011:00005",
  "USGS:05082500:00011:00025",
  "USGS:05082500:00011:00027",
  "USGS:05082500:00011:00028",
  "USGS:05082500:00011:00029",
  "USGS:05082625:00011:00002",
  "USGS:05082625:00011:00005",
  "USGS:05082625:00011:00018",
  "USGS:05084000:00011:00001",
  "USGS:05084000:00011:00003",
  "USGS:05085000:00011:00001",
  "USGS:05085000:00011:00003",
  "USGS:05090000:00011:00001",
  "USGS:05090000:00011:00004",
  "USGS:05090000:00011:00005",
  "USGS:05092000:00011:00003",
  "USGS:05092000:00011:00006",
  "USGS:05099400:00011:00001",
  "USGS:05099400:00011:00002",
  "USGS:05099400:00011:00016",
  "USGS:05099600:00011:00002",
  "USGS:05099600:00011:00003",
  "USGS:05099600:00011:00015",
  "USGS:05100000:00011:00001",
  "USGS:05100000:00011:00004",
  "USGS:05100000:00011:00007",
  "USGS:05101000:00011:00001",
  "USGS:05101000:00011:00003",
  "USGS:05102490:00011:00001",
  "USGS:05113600:00011:00001",
  "USGS:05113600:00011:00003",
  "USGS:05113750:00011:00004",
  "USGS:05114000:00011:00002",
  "USGS:05114000:00011:00008",
  "USGS:05115500:00011:00001",
  "USGS:05116000:00011:00002",
  "USGS:05116000:00011:00005",
  "USGS:05116500:00011:00001",
  "USGS:05116500:00011:00004",
  "USGS:05117500:00011:00001",
  "USGS:05117500:00011:00003",
  "USGS:05120000:00011:00002",
  "USGS:05120000:00011:00006",
  "USGS:05120500:00011:00001",
  "USGS:05120500:00011:00003",
  "USGS:05122000:00011:00001",
  "USGS:05122000:00011:00007",
  "USGS:05123400:00011:00001",
  "USGS:05123400:00011:00007",
  "USGS:05123510:00011:00002",
  "USGS:05123510:00011:00005",
  "USGS:05124000:00011:00002",
  "USGS:05124000:00011:00007",
  "USGS:06329595:00011:00001",
  "USGS:06329595:00011:00002",
  "USGS:06329597:00011:00002",
  "USGS:06329597:00011:00001",
  "USGS:06329597:00011:00014",
  "USGS:06329597:00011:00003",
  "USGS:06329610:00011:00002",
  "USGS:06330000:00011:00001",
  "USGS:06330000:00011:00003",
  "USGS:06330110:00011:00002",
  "USGS:06331000:00011:00001",
  "USGS:06331000:00011:00014",
  "USGS:06332000:00011:00002",
  "USGS:06332000:00011:00004",
  "USGS:06332515:00011:00002",
  "USGS:06332515:00011:00006",
  "USGS:06335500:00011:00002",
  "USGS:06335500:00011:00006",
  "USGS:06335750:00011:00001",
  "USGS:06335750:00011:00003",
  "USGS:06336000:00011:00001",
  "USGS:06336000:00011:00002",
  "USGS:06336000:00011:00005",
  "USGS:06336000:00011:00019",
  "USGS:06336000:00011:00020",
  "USGS:06336000:00011:00021",
  "USGS:06336600:00011:00001",
  "USGS:06336600:00011:00003",
  "USGS:03028500:00011:00017",
  "USGS:03028500:00011:00004",
  "USGS:03028500:00011:00003",
  "USGS:01155500:00011:00001",
  "USGS:01155500:00011:00003",
  "USGS:01155910:00011:00002",
  "USGS:01155910:00011:00005",
  "USGS:01334000:00011:00001",
  "USGS:01334000:00011:00003",
  "USGS:021720698:00011:00003",
  "USGS:021720698:00011:00004",
  "USGS:021720698:00011:00001",
  "USGS:021720698:00011:00002",
  "USGS:04279490:00011:00001",
  "USGS:04280000:00011:00001",
  "USGS:04280000:00011:00004",
  "USGS:04282000:00011:00001",
  "USGS:04282000:00011:00003",
  "USGS:04282500:00011:00001",
  "USGS:04282500:00011:00003",
  "USGS:04282525:00011:00003",
  "USGS:04282525:00011:00002",
  "USGS:04282525:00011:00004",
  "USGS:04282650:00011:00002",
  "USGS:04282650:00011:00001",
  "USGS:0505152130:00011:00003",
  "USGS:0505152130:00011:00001",
  "USGS:05051522:00011:00002",
  "USGS:05051522:00011:00001",
  "USGS:05051600:00011:00001",
  "USGS:05051600:00011:00003",
  "USGS:05052000:00011:00001" ;

 v00065_description =
  "USGS:02339495:00011:00002",
  "USGS:02339495:00011:00001",
  "USGS:02342500:00011:00001",
  "USGS:02342500:00011:00002",
  "USGS:0234296910:00011:00002",
  "USGS:023432415:00011:00016",
  "USGS:023432415:00011:00003",
  "USGS:023432415:00011:00002",
  "USGS:023432415:00011:00001",
  "USGS:023432415:00011:00017",
  "USGS:023432415:00011:00018",
  "USGS:02361000:00011:00010",
  "USGS:02361000:00011:00011",
  "USGS:02361000:00011:00002",
  "USGS:02361000:00011:00003",
  "USGS:02361500:00011:00005",
  "USGS:02361500:00011:00006",
  "USGS:02361500:00011:00001",
  "USGS:02361500:00011:00002",
  "USGS:02362000:00011:00002",
  "USGS:02362240:00011:00001",
  "USGS:02362240:00011:00002",
  "USGS:02363000:00011:00001",
  "USGS:02363000:00011:00002",
  "USGS:02364000:00011:00001",
  "USGS:02364500:00011:00005",
  "USGS:02364500:00011:00006",
  "USGS:02364500:00011:00001",
  "USGS:02364500:00011:00002",
  "USGS:02369800:00011:00002",
  "USGS:02369800:00011:00003",
  "USGS:02371500:00011:00005",
  "USGS:02371500:00011:00006",
  "USGS:02372250:00011:00001",
  "USGS:02372250:00011:00002",
  "USGS:02372422:00011:00005",
  "USGS:02372422:00011:00004",
  "USGS:02372430:00011:00003",
  "USGS:02372430:00011:00001",
  "USGS:02373000:00011:00001",
  "USGS:02373000:00011:00002",
  "USGS:02374250:00011:00002",
  "USGS:02374250:00011:00001",
  "USGS:02374500:00011:00001",
  "USGS:02374500:00011:00002",
  "USGS:02374700:00011:00004",
  "USGS:02374700:00011:00002",
  "USGS:02374700:00011:00001",
  "USGS:02374745:00011:00002",
  "USGS:02374745:00011:00001",
  "USGS:02374950:00011:00002",
  "USGS:02374950:00011:00001",
  "USGS:02376500:00011:00002",
  "USGS:02376500:00011:00001",
  "USGS:02377560:00011:00001",
  "USGS:02377570:00011:00002",
  "USGS:02377570:00011:00001",
  "USGS:02377750:00011:00001",
  "USGS:02378170:00011:00002",
  "USGS:02378170:00011:00001",
  "USGS:02378300:00011:00002",
  "USGS:02378300:00011:00001",
  "USGS:02378500:00011:00003",
  "USGS:02378500:00011:00001",
  "USGS:02378500:00011:00002",
  "USGS:02397530:00011:00001",
  "USGS:02397530:00011:00007",
  "USGS:02397530:00011:00026",
  "USGS:02397530:00011:00027",
  "USGS:02397530:00011:00017",
  "USGS:02397530:00011:00002",
  "USGS:02397530:00011:00003",
  "USGS:02397530:00011:00004",
  "USGS:02398300:00011:00001",
  "USGS:02398300:00011:00002",
  "USGS:02399200:00011:00001",
  "USGS:02399200:00011:00002",
  "USGS:02399500:00011:00002",
  "USGS:02400100:00011:00001",
  "USGS:02400100:00011:00002",
  "USGS:02400496:00011:00002",
  "USGS:02400500:00011:00003",
  "USGS:02400680:00011:00002",
  "USGS:02400680:00011:00001",
  "USGS:02401000:00011:00001",
  "USGS:02401000:00011:00002",
  "USGS:02401390:00011:00001",
  "USGS:02401390:00011:00002",
  "USGS:02401895:00011:00002",
  "USGS:02401895:00011:00001",
  "USGS:02403310:00011:00001",
  "USGS:07176321:00011:00002",
  "USGS:02404400:00011:00001",
  "USGS:02404400:00011:00002",
  "USGS:02405500:00011:00004",
  "USGS:02405500:00011:00001",
  "USGS:02405500:00011:00002",
  "USGS:02406500:00011:00001",
  "USGS:02406500:00011:00002",
  "USGS:02406930:00011:00002",
  "USGS:02406930:00011:00001",
  "USGS:02407000:00011:00004",
  "USGS:02407000:00011:00002",
  "USGS:02407000:00011:00003",
  "USGS:02407514:00011:00004",
  "USGS:02407514:00011:00002",
  "USGS:02407514:00011:00001",
  "USGS:02407526:00011:00001",
  "USGS:02408150:00011:00001",
  "USGS:02408540:00011:00001",
  "USGS:02408540:00011:00002",
  "USGS:01118300:00011:00004",
  "USGS:01118300:00011:00016",
  "USGS:01118300:00011:00001",
  "USGS:01118300:00011:00003",
  "USGS:01119382:00011:00013",
  "USGS:01119382:00011:00015",
  "USGS:01119382:00011:00009",
  "USGS:01119382:00011:00002",
  "USGS:01119382:00011:00001",
  "USGS:01119500:00011:00002",
  "USGS:01119500:00011:00005",
  "USGS:01120790:00011:00004",
  "USGS:01120790:00011:00005",
  "USGS:01120790:00011:00007",
  "USGS:01120790:00011:00001",
  "USGS:01120790:00011:00002",
  "USGS:01121000:00011:00001",
  "USGS:01121000:00011:00003",
  "USGS:01121330:00011:00001",
  "USGS:01121330:00011:00002",
  "USGS:01121500:00011:00002",
  "USGS:02471078:00011:00002",
  "USGS:02471078:00011:00001",
  "USGS:02479945:00011:00002",
  "USGS:02479945:00011:00001",
  "USGS:02479980:00011:00002",
  "USGS:02479980:00011:00001",
  "USGS:02480002:00011:00002",
  "USGS:02480002:00011:00001",
  "USGS:03572690:00011:00002",
  "USGS:03572690:00011:00001",
  "USGS:03574500:00011:00004",
  "USGS:03574500:00011:00005",
  "USGS:0357479650:00011:00001",
  "USGS:03575100:00011:00002",
  "USGS:03575100:00011:00001",
  "USGS:0357526200:00011:00003",
  "USGS:0357526200:00011:00002",
  "USGS:0357526200:00011:00001",
  "USGS:03575272:00011:00004",
  "USGS:03575272:00011:00002",
  "USGS:03575272:00011:00001",
  "USGS:03575500:00011:00002",
  "USGS:0357568650:00011:00003",
  "USGS:0357568650:00011:00002",
  "USGS:0357568650:00011:00001",
  "USGS:0357568980:00011:00003",
  "USGS:0357568980:00011:00002",
  "USGS:0357568980:00011:00001",
  "USGS:03575700:00011:00001",
  "USGS:03575700:00011:00002",
  "USGS:03575700:00011:00003",
  "USGS:03575830:00011:00001",
  "USGS:03575830:00011:00002",
  "USGS:03575830:00011:00003",
  "USGS:0357586650:00011:00003",
  "USGS:0357586650:00011:00002",
  "USGS:0357586650:00011:00001",
  "USGS:0357587090:00011:00003",
  "USGS:0357587090:00011:00002",
  "USGS:0357587090:00011:00001",
  "USGS:0357587140:00011:00003",
  "USGS:0357587140:00011:00002",
  "USGS:0357587140:00011:00001",
  "USGS:0357587400:00011:00003",
  "USGS:0357587400:00011:00002",
  "USGS:0357587400:00011:00001",
  "USGS:0357587728:00011:00001",
  "USGS:0357587728:00011:00002",
  "USGS:0357587728:00011:00003",
  "USGS:02411600:00011:00003",
  "USGS:03575890:00011:00001",
  "USGS:03575890:00011:00002",
  "USGS:03575890:00011:00003",
  "USGS:0357591500:00011:00003",
  "USGS:0357591500:00011:00002",
  "USGS:0357591500:00011:00001",
  "USGS:03575950:00011:00001",
  "USGS:03575950:00011:00002",
  "USGS:03575950:00011:00003",
  "USGS:03575980:00011:00001",
  "USGS:03575980:00011:00003",
  "USGS:03575980:00011:00002",
  "USGS:03576250:00011:00001",
  "USGS:03576250:00011:00002",
  "USGS:03576500:00011:00002",
  "USGS:03576500:00011:00003",
  "USGS:03577150:00011:00002",
  "USGS:03577225:00011:00002",
  "USGS:03577225:00011:00001",
  "USGS:03586500:00011:00002",
  "USGS:03586500:00011:00003",
  "USGS:03589500:00011:00003",
  "USGS:03590000:00011:00002",
  "USGS:03592500:00011:00003",
  "USGS:322047086214301:00011:00001",
  "USGS:322500085551201:00011:00001",
  "USGS:332934086353801:00011:00001",
  "USGS:333103086524501:00011:00001",
  "USGS:333204087324601:00011:00001",
  "USGS:333205086493701:00011:00002",
  "USGS:333437086430801:00011:00001",
  "USGS:335929087021001:00011:00001",
  "USGS:340618086344001:00011:00001",
  "USGS:342718087285601:00011:00001",
  "USGS:343843085403201:00011:00001",
  "USGS:02204520:00011:00015",
  "USGS:02204520:00011:00005",
  "USGS:02204520:00011:00016",
  "USGS:02204520:00011:00017",
  "USGS:02204520:00011:00002",
  "USGS:02204520:00011:00001",
  "USGS:02205000:00011:00006",
  "USGS:02205865:00011:00004",
  "USGS:02205865:00011:00003",
  "USGS:02205865:00011:00002",
  "USGS:02205865:00011:00001",
  "USGS:02205865:00011:00005",
  "USGS:02207120:00011:00006",
  "USGS:02207120:00011:00003",
  "USGS:02207120:00011:00002",
  "USGS:02207120:00011:00001",
  "USGS:02207120:00011:00007",
  "USGS:02207130:00011:00005",
  "USGS:02207130:00011:00004",
  "USGS:02207135:00011:00007",
  "USGS:02207135:00011:00005",
  "USGS:02207135:00011:00004",
  "USGS:02207135:00011:00008",
  "USGS:02207135:00011:00009",
  "USGS:02412000:00011:00001",
  "USGS:02412000:00011:00002",
  "USGS:02413300:00011:00001",
  "USGS:02413300:00011:00002",
  "USGS:02414500:00011:00001",
  "USGS:02414500:00011:00002",
  "USGS:02414715:00011:00001",
  "USGS:02414715:00011:00002",
  "USGS:02415000:00011:00001",
  "USGS:02415000:00011:00002",
  "USGS:02418230:00011:00002",
  "USGS:02418230:00011:00001",
  "USGS:02418760:00011:00002",
  "USGS:02418760:00011:00001",
  "USGS:02419000:00011:00001",
  "USGS:02419000:00011:00002",
  "USGS:02419500:00011:00002",
  "USGS:02419890:00011:00004",
  "USGS:02419890:00011:00002",
  "USGS:02419890:00011:00001",
  "USGS:02419890:00011:00006",
  "USGS:02419890:00011:00008",
  "USGS:02419988:00011:00001",
  "USGS:02420000:00011:00007",
  "USGS:02420000:00011:00003",
  "USGS:02420000:00011:00004",
  "USGS:02420490:00011:00001",
  "USGS:02421000:00011:00001",
  "USGS:02421000:00011:00002",
  "USGS:02421350:00011:00002",
  "USGS:02421350:00011:00001",
  "USGS:02421351:00011:00002",
  "USGS:02422500:00011:00001",
  "USGS:02422500:00011:00002",
  "USGS:02423000:00011:00003",
  "USGS:02423110:00011:00001",
  "USGS:02423110:00011:00003",
  "USGS:02423130:00011:00003",
  "USGS:02423130:00011:00002",
  "USGS:02423130:00011:00001",
  "USGS:02423130:00011:00004",
  "USGS:02423130:00011:00005",
  "USGS:02423160:00011:00003",
  "USGS:02423160:00011:00002",
  "USGS:02423160:00011:00001",
  "USGS:02423160:00011:00004",
  "USGS:02423160:00011:00005",
  "USGS:02423380:00011:00006",
  "USGS:02423380:00011:00007",
  "USGS:02423397:00011:00004",
  "USGS:02423397:00011:00002",
  "USGS:02423397:00011:00001",
  "USGS:02423397:00011:00005",
  "USGS:02423397:00011:00006",
  "USGS:02423400:00011:00004",
  "USGS:02423400:00011:00002",
  "USGS:02423414:00011:00002",
  "USGS:02423414:00011:00001",
  "USGS:02423425:00011:00002",
  "USGS:02423425:00011:00001",
  "USGS:07176321:00011:00001",
  "USGS:02423496:00011:00003",
  "USGS:02423496:00011:00002",
  "USGS:02423496:00011:00001",
  "USGS:02423496:00011:00004",
  "USGS:02423496:00011:00005",
  "USGS:02423500:00011:00001",
  "USGS:02423500:00011:00002",
  "USGS:0242354750:00011:00002",
  "USGS:0242354750:00011:00001",
  "USGS:02423555:00011:00002",
  "USGS:02423555:00011:00001",
  "USGS:02423630:00011:00001",
  "USGS:02423630:00011:00002",
  "USGS:02424000:00011:00004",
  "USGS:02424000:00011:00005",
  "USGS:02424590:00011:00001",
  "USGS:02425000:00011:00001",
  "USGS:02425000:00011:00002",
  "USGS:02427250:00011:00002",
  "USGS:02427250:00011:00001",
  "USGS:02427505:00011:00002",
  "USGS:02427505:00011:00001",
  "USGS:02427506:00011:00002",
  "USGS:02427830:00011:00002",
  "USGS:02427830:00011:00001",
  "USGS:02428400:00011:00002",
  "USGS:02428400:00011:00003",
  "USGS:02428400:00011:00006",
  "USGS:02428400:00011:00007",
  "USGS:02428400:00011:00008",
  "USGS:02428400:00011:00009",
  "USGS:02428400:00011:00010",
  "USGS:02428400:00011:00011",
  "USGS:02428401:00011:00002",
  "USGS:02438000:00011:00001",
  "USGS:02438000:00011:00002",
  "USGS:02444160:00011:00001",
  "USGS:02444160:00011:00003",
  "USGS:02444160:00011:00005",
  "USGS:02444160:00011:00006",
  "USGS:02444160:00011:00007",
  "USGS:02444160:00011:00008",
  "USGS:02444161:00011:00001",
  "USGS:02446500:00011:00001",
  "USGS:02446500:00011:00002",
  "USGS:02447025:00011:00001",
  "USGS:02447025:00011:00003",
  "USGS:02447025:00011:00005",
  "USGS:02447025:00011:00006",
  "USGS:02447025:00011:00007",
  "USGS:02447025:00011:00008",
  "USGS:02447025:00011:00009",
  "USGS:02447026:00011:00001",
  "USGS:02448500:00011:00001",
  "USGS:02448500:00011:00002",
  "USGS:02448900:00011:00002",
  "USGS:02448900:00011:00001",
  "USGS:02449882:00011:00002",
  "USGS:02449882:00011:00001",
  "USGS:02193340:00011:00001",
  "USGS:02193340:00011:00002",
  "USGS:15085100:00011:00007",
  "USGS:15085100:00011:00002",
  "USGS:15085100:00011:00005",
  "USGS:15099900:00011:00013",
  "USGS:15099900:00011:00015",
  "USGS:15099900:00011:00001",
  "USGS:15099900:00011:00002",
  "USGS:15099900:00011:00003",
  "USGS:15100000:00011:00012",
  "USGS:15100000:00011:00001",
  "USGS:15100000:00011:00002",
  "USGS:15100000:00011:00003",
  "USGS:15101490:00011:00002",
  "USGS:15101490:00011:00003",
  "USGS:15129120:00011:00005",
  "USGS:15129120:00011:00015",
  "USGS:15129120:00011:00016",
  "USGS:15129120:00011:00003",
  "USGS:15129120:00011:00001",
  "USGS:15129120:00011:00002",
  "USGS:15129120:00011:00006",
  "USGS:15129500:00011:00008",
  "USGS:15129500:00011:00002",
  "USGS:15129500:00011:00019",
  "USGS:15129500:00011:00004",
  "USGS:15129500:00011:00006",
  "USGS:15129500:00011:00009",
  "USGS:15200280:00011:00001",
  "USGS:15200280:00011:00002",
  "USGS:15200280:00011:00003",
  "USGS:15214000:00011:00016",
  "USGS:15214000:00011:00017",
  "USGS:15214000:00011:00020",
  "USGS:15214000:00011:00005",
  "USGS:15214000:00011:00002",
  "USGS:15214000:00011:00003",
  "USGS:15225997:00011:00001",
  "USGS:15225997:00011:00002",
  "USGS:15225997:00011:00005",
  "USGS:15226620:00011:00002",
  "USGS:15226620:00011:00001",
  "USGS:15236895:00011:00002",
  "USGS:15236895:00011:00004",
  "USGS:15236895:00011:00025",
  "USGS:15236895:00011:00014",
  "USGS:15236895:00011:00016",
  "USGS:15236895:00011:00020",
  "USGS:15236895:00011:00026",
  "USGS:15236895:00011:00019",
  "USGS:15236895:00011:00001",
  "USGS:15236895:00011:00023",
  "USGS:15236900:00011:00005",
  "USGS:15236900:00011:00016",
  "USGS:15236900:00011:00001",
  "USGS:15236900:00011:00003",
  "USGS:15237730:00011:00003",
  "USGS:15237730:00011:00014",
  "USGS:15237730:00011:00001",
  "USGS:15238648:00011:00003",
  "USGS:15238648:00011:00004",
  "USGS:15238648:00011:00001",
  "USGS:15238648:00011:00002",
  "USGS:15238648:00011:00008",
  "USGS:15238990:00011:00004",
  "USGS:15238990:00011:00002",
  "USGS:15238990:00011:00007",
  "USGS:15238990:00011:00009",
  "USGS:15239001:00011:00004",
  "USGS:15239001:00011:00020",
  "USGS:15239001:00011:00021",
  "USGS:15239001:00011:00019",
  "USGS:15239001:00011:00005",
  "USGS:15239001:00011:00018",
  "USGS:15239001:00011:00002",
  "USGS:15239001:00011:00001",
  "USGS:15239001:00011:00017",
  "USGS:15239001:00011:00007",
  "USGS:15239050:00011:00005",
  "USGS:15239050:00011:00001",
  "USGS:15239050:00011:00002",
  "USGS:15239050:00011:00008",
  "USGS:15239060:00011:00004",
  "USGS:15239060:00011:00002",
  "USGS:15239060:00011:00001",
  "USGS:15239060:00011:00007",
  "USGS:15239070:00011:00002",
  "USGS:15239070:00011:00007",
  "USGS:15239070:00011:00003",
  "USGS:15239070:00011:00005",
  "USGS:15239070:00011:00014",
  "USGS:15239070:00011:00006",
  "USGS:15239900:00011:00004",
  "USGS:15239900:00011:00002",
  "USGS:15243900:00011:00005",
  "USGS:15243900:00011:00001",
  "USGS:15243900:00011:00003",
  "USGS:15258000:00011:00003",
  "USGS:15258000:00011:00017",
  "USGS:15258000:00011:00006",
  "USGS:15258000:00011:00004",
  "USGS:15258000:00011:00002",
  "USGS:15261000:00011:00003",
  "USGS:15261000:00011:00001",
  "USGS:15261000:00011:00002",
  "USGS:15266110:00011:00003",
  "USGS:15266110:00011:00002",
  "USGS:15266110:00011:00001",
  "USGS:15266300:00011:00017",
  "USGS:15266300:00011:00023",
  "USGS:15266300:00011:00001",
  "USGS:15266300:00011:00005",
  "USGS:15271000:00011:00015",
  "USGS:15271000:00011:00004",
  "USGS:15271000:00011:00005",
  "USGS:15274600:00011:00006",
  "USGS:15274600:00011:00005",
  "USGS:15275100:00011:00010",
  "USGS:15275100:00011:00007",
  "USGS:15276000:00011:00008",
  "USGS:15276000:00011:00002",
  "USGS:15276000:00011:00004",
  "USGS:15278000:00011:00002",
  "USGS:15278000:00011:00001",
  "USGS:15283700:00011:00014",
  "USGS:15283700:00011:00001",
  "USGS:15283700:00011:00002",
  "USGS:15284000:00011:00001",
  "USGS:15284000:00011:00002",
  "USGS:15284000:00011:00006",
  "USGS:15290000:00011:00003",
  "USGS:15290000:00011:00014",
  "USGS:15291700:00011:00012",
  "USGS:15291700:00011:00017",
  "USGS:15291700:00011:00001",
  "USGS:15291700:00011:00002",
  "USGS:15292000:00011:00005",
  "USGS:15292000:00011:00020",
  "USGS:15292000:00011:00001",
  "USGS:15292400:00011:00001",
  "USGS:15292400:00011:00002",
  "USGS:15292400:00011:00003",
  "USGS:15292400:00011:00013",
  "USGS:15292700:00011:00001",
  "USGS:15292700:00011:00019",
  "USGS:15292700:00011:00008",
  "USGS:15292700:00011:00002",
  "USGS:15292700:00011:00003",
  "USGS:15292700:00011:00020",
  "USGS:15292780:00011:00004",
  "USGS:15292780:00011:00005",
  "USGS:15292780:00011:00006",
  "USGS:15292780:00011:00015",
  "USGS:15292780:00011:00003",
  "USGS:15292800:00011:00016",
  "USGS:15292800:00011:00003",
  "USGS:15292800:00011:00006",
  "USGS:15292800:00011:00001",
  "USGS:15293200:00011:00013",
  "USGS:15293200:00011:00014",
  "USGS:15293200:00011:00003",
  "USGS:15293200:00011:00001",
  "USGS:15293200:00011:00002",
  "USGS:15293700:00011:00003",
  "USGS:15293700:00011:00001",
  "USGS:15293700:00011:00002",
  "USGS:15294005:00011:00017",
  "USGS:15294005:00011:00003",
  "USGS:15294005:00011:00006",
  "USGS:15294005:00011:00002",
  "USGS:15295700:00011:00004",
  "USGS:15295700:00011:00022",
  "USGS:15295700:00011:00018",
  "USGS:15295700:00011:00015",
  "USGS:15295700:00011:00016",
  "USGS:15297610:00011:00003",
  "USGS:15297610:00011:00001",
  "USGS:15297610:00011:00002",
  "USGS:15298040:00011:00001",
  "USGS:15298040:00011:00019",
  "USGS:15298040:00011:00002",
  "USGS:15298040:00011:00003",
  "USGS:15298040:00011:00017",
  "USGS:15300100:00011:00003",
  "USGS:15300100:00011:00013",
  "USGS:15300100:00011:00001",
  "USGS:15300100:00011:00002",
  "USGS:15300250:00011:00014",
  "USGS:15300250:00011:00016",
  "USGS:15300250:00011:00003",
  "USGS:15300250:00011:00001",
  "USGS:15300250:00011:00013",
  "USGS:15300300:00011:00014",
  "USGS:15300300:00011:00016",
  "USGS:15300300:00011:00012",
  "USGS:15300300:00011:00002",
  "USGS:15300300:00011:00013",
  "USGS:15302000:00011:00016",
  "USGS:15302000:00011:00018",
  "USGS:15302000:00011:00014",
  "USGS:15302000:00011:00004",
  "USGS:15302000:00011:00005",
  "USGS:01096000:00011:00001",
  "USGS:01096000:00011:00003",
  "USGS:01122000:00011:00001",
  "USGS:01122000:00011:00005",
  "USGS:01122500:00011:00001",
  "USGS:01122500:00011:00003",
  "USGS:01123000:00011:00001",
  "USGS:01123000:00011:00003",
  "USGS:011230695:00011:00002",
  "USGS:011230695:00011:00014",
  "USGS:01124000:00011:00001",
  "USGS:01124000:00011:00003",
  "USGS:01124151:00011:00014",
  "USGS:01124151:00011:00013",
  "USGS:01124151:00011:00001",
  "USGS:01124151:00011:00005",
  "USGS:01125100:00011:00002",
  "USGS:01125100:00011:00001",
  "USGS:01125490:00011:00001",
  "USGS:01125490:00011:00002",
  "USGS:01125500:00011:00004",
  "USGS:01125500:00011:00005",
  "USGS:01127000:00011:00002",
  "USGS:01127000:00011:00005",
  "USGS:01127500:00011:00016",
  "USGS:01127500:00011:00001",
  "USGS:01127500:00011:00006",
  "USGS:011277905:00011:00002",
  "USGS:011277905:00011:00001",
  "USGS:01184000:00011:00002",
  "USGS:01184000:00011:00005",
  "USGS:01184100:00011:00017",
  "USGS:01184100:00011:00019",
  "USGS:01184100:00011:00001",
  "USGS:01184100:00011:00007",
  "USGS:01184490:00011:00001",
  "USGS:01184490:00011:00004",
  "USGS:01186000:00011:00002",
  "USGS:01186000:00011:00005",
  "USGS:01186500:00011:00001",
  "USGS:01186500:00011:00004",
  "USGS:01187300:00011:00005",
  "USGS:01187300:00011:00006",
  "USGS:01187300:00011:00001",
  "USGS:01187300:00011:00002",
  "USGS:01188000:00011:00002",
  "USGS:01188000:00011:00004",
  "USGS:01188090:00011:00002",
  "USGS:01188090:00011:00003",
  "USGS:01189213:00011:00001",
  "USGS:01189995:00011:00002",
  "USGS:01189995:00011:00005",
  "USGS:01190070:00011:00005",
  "USGS:01191000:00011:00001",
  "USGS:01191000:00011:00002",
  "USGS:01192500:00011:00002",
  "USGS:01192500:00011:00014",
  "USGS:01192883:00011:00016",
  "USGS:01192883:00011:00018",
  "USGS:01192883:00011:00001",
  "USGS:01192883:00011:00006",
  "USGS:01193050:00011:00006",
  "USGS:01193050:00011:00026",
  "USGS:01193050:00011:00035",
  "USGS:01193050:00011:00012",
  "USGS:01193050:00011:00011",
  "USGS:01193050:00011:00009",
  "USGS:01193050:00011:00007",
  "USGS:01193050:00011:00010",
  "USGS:01193050:00011:00038",
  "USGS:01193050:00011:00037",
  "USGS:01193050:00011:00041",
  "USGS:01193500:00011:00001",
  "USGS:01193500:00011:00011",
  "USGS:01193500:00011:00002",
  "USGS:01193500:00011:00003",
  "USGS:01194000:00011:00005",
  "USGS:01194000:00011:00004",
  "USGS:01194000:00011:00001",
  "USGS:01194000:00011:00002",
  "USGS:01194500:00011:00017",
  "USGS:01194500:00011:00016",
  "USGS:01194500:00011:00003",
  "USGS:01194500:00011:00001",
  "USGS:01194500:00011:00002",
  "USGS:01194750:00011:00003",
  "USGS:01194750:00011:00010",
  "USGS:01194750:00011:00013",
  "USGS:01194750:00011:00001",
  "USGS:01194750:00011:00004",
  "USGS:01194750:00011:00011",
  "USGS:01194750:00011:00014",
  "USGS:01194750:00011:00006",
  "USGS:01194750:00011:00007",
  "USGS:01194750:00011:00008",
  "USGS:01194750:00011:00009",
  "USGS:01194750:00011:00005",
  "USGS:01194750:00011:00012",
  "USGS:01194750:00011:00015",
  "USGS:01194796:00011:00004",
  "USGS:01194796:00011:00006",
  "USGS:01194796:00011:00001",
  "USGS:01194796:00011:00005",
  "USGS:01194796:00011:00007",
  "USGS:01194796:00011:00009",
  "USGS:01194796:00011:00010",
  "USGS:01195100:00011:00004",
  "USGS:01195100:00011:00001",
  "USGS:01195100:00011:00003",
  "USGS:01195490:00011:00011",
  "USGS:01195490:00011:00002",
  "USGS:01195490:00011:00003",
  "USGS:01196500:00011:00001",
  "USGS:01196500:00011:00017",
  "USGS:01196500:00011:00014",
  "USGS:01196500:00011:00002",
  "USGS:01196500:00011:00003",
  "USGS:01196500:00011:00004",
  "USGS:01196500:00011:00016",
  "USGS:01196561:00011:00002",
  "USGS:01196561:00011:00001",
  "USGS:01196620:00011:00001",
  "USGS:01196620:00011:00003",
  "USGS:01199000:00011:00019",
  "USGS:01199000:00011:00018",
  "USGS:01199000:00011:00002",
  "USGS:01199000:00011:00003",
  "USGS:01199050:00011:00001",
  "USGS:01199050:00011:00003",
  "USGS:01200500:00011:00002",
  "USGS:01200500:00011:00008",
  "USGS:02457595:00011:00005",
  "USGS:01200600:00011:00002",
  "USGS:01200600:00011:00009",
  "USGS:01200600:00011:00003",
  "USGS:01200600:00011:00011",
  "USGS:01201487:00011:00014",
  "USGS:01201487:00011:00017",
  "USGS:01201487:00011:00003",
  "USGS:01201487:00011:00002",
  "USGS:01201487:00011:00001",
  "USGS:01201487:00011:00015",
  "USGS:01201487:00011:00016",
  "USGS:01202501:00011:00014",
  "USGS:01202501:00011:00002",
  "USGS:01202501:00011:00001",
  "USGS:012035055:00011:00002",
  "USGS:012035055:00011:00001",
  "USGS:01203510:00011:00001",
  "USGS:01203510:00011:00002",
  "USGS:01203600:00011:00001",
  "USGS:01203600:00011:00003",
  "USGS:01203805:00011:00019",
  "USGS:01203805:00011:00018",
  "USGS:01203805:00011:00001",
  "USGS:01203805:00011:00003",
  "USGS:01204000:00011:00002",
  "USGS:01204000:00011:00005",
  "USGS:07294800:00011:00001",
  "USGS:02450000:00011:00002",
  "USGS:02450000:00011:00003",
  "USGS:02450180:00011:00002",
  "USGS:02450180:00011:00003",
  "USGS:02450250:00011:00006",
  "USGS:02450250:00011:00001",
  "USGS:02450250:00011:00002",
  "USGS:02450825:00011:00002",
  "USGS:02450825:00011:00003",
  "USGS:02453000:00011:00003",
  "USGS:02453000:00011:00004",
  "USGS:02453500:00011:00009",
  "USGS:02453500:00011:00001",
  "USGS:02453500:00011:00002",
  "USGS:02454055:00011:00002",
  "USGS:02454055:00011:00001",
  "USGS:02455000:00011:00002",
  "USGS:02455000:00011:00003",
  "USGS:02455185:00011:00002",
  "USGS:02455185:00011:00001",
  "USGS:02455980:00011:00003",
  "USGS:02455980:00011:00001",
  "USGS:02455980:00011:00002",
  "USGS:02455980:00011:00004",
  "USGS:02455980:00011:00005",
  "USGS:02456500:00011:00002",
  "USGS:02456500:00011:00003",
  "USGS:02457000:00011:00002",
  "USGS:02457000:00011:00003",
  "USGS:02457595:00011:00003",
  "USGS:02457595:00011:00002",
  "USGS:02457595:00011:00001",
  "USGS:02457595:00011:00004",
  "USGS:02458148:00011:00004",
  "USGS:02458148:00011:00002",
  "USGS:02458148:00011:00001",
  "USGS:02458148:00011:00005",
  "USGS:02458190:00011:00002",
  "USGS:02458190:00011:00001",
  "USGS:02458300:00011:00003",
  "USGS:02458300:00011:00002",
  "USGS:02458450:00011:00004",
  "USGS:02458450:00011:00002",
  "USGS:02458450:00011:00003",
  "USGS:02458450:00011:00005",
  "USGS:02458450:00011:00006",
  "USGS:02458502:00011:00004",
  "USGS:02458502:00011:00002",
  "USGS:02458502:00011:00001",
  "USGS:02458502:00011:00005",
  "USGS:02458600:00011:00002",
  "USGS:02458600:00011:00001",
  "USGS:02461500:00011:00002",
  "USGS:02461500:00011:00003",
  "USGS:02462000:00011:00002",
  "USGS:02462000:00011:00003",
  "USGS:02462500:00011:00008",
  "USGS:02462500:00011:00003",
  "USGS:02462501:00011:00001",
  "USGS:02462951:00011:00005",
  "USGS:02462951:00011:00004",
  "USGS:02462952:00011:00001",
  "USGS:02464000:00011:00002",
  "USGS:02464000:00011:00003",
  "USGS:02464146:00011:00002",
  "USGS:02464146:00011:00001",
  "USGS:02464360:00011:00002",
  "USGS:02464360:00011:00003",
  "USGS:02464660:00011:00002",
  "USGS:02464660:00011:00001",
  "USGS:02464800:00011:00011",
  "USGS:02464800:00011:00003",
  "USGS:02464800:00011:00007",
  "USGS:02465000:00011:00003",
  "USGS:02465000:00011:00004",
  "USGS:02465005:00011:00001",
  "USGS:02465292:00011:00002",
  "USGS:02465292:00011:00001",
  "USGS:02465493:00011:00001",
  "USGS:02465493:00011:00002",
  "USGS:02466030:00011:00001",
  "USGS:02466030:00011:00003",
  "USGS:02466030:00011:00005",
  "USGS:02466030:00011:00006",
  "USGS:02466030:00011:00007",
  "USGS:02466030:00011:00008",
  "USGS:02466030:00011:00009",
  "USGS:02466030:00011:00010",
  "USGS:02466031:00011:00003",
  "USGS:02467000:00011:00001",
  "USGS:02467000:00011:00002",
  "USGS:02467001:00011:00002",
  "USGS:02467500:00011:00001",
  "USGS:02467500:00011:00002",
  "USGS:02469525:00011:00004",
  "USGS:02469525:00011:00001",
  "USGS:02469761:00011:00001",
  "USGS:02469761:00011:00002",
  "USGS:02469761:00011:00005",
  "USGS:02469761:00011:00006",
  "USGS:02469761:00011:00007",
  "USGS:02469761:00011:00008",
  "USGS:02469761:00011:00009",
  "USGS:02469761:00011:00010",
  "USGS:02469761:00011:00011",
  "USGS:02469761:00011:00012",
  "USGS:02469762:00011:00002",
  "USGS:02469800:00011:00001",
  "USGS:02469800:00011:00002",
  "USGS:02470050:00011:00001",
  "USGS:02470072:00011:00003",
  "USGS:02470072:00011:00002",
  "USGS:02470629:00011:00005",
  "USGS:02470629:00011:00004",
  "USGS:02470629:00011:00003",
  "USGS:02470629:00011:00026",
  "USGS:02470630:00011:00001",
  "USGS:02471001:00011:00001",
  "USGS:02471001:00011:00002",
  "USGS:02471019:00011:00002",
  "USGS:02471019:00011:00004",
  "USGS:03613000:00011:00003",
  "USGS:03613000:00011:00001",
  "USGS:01205500:00011:00002",
  "USGS:01205500:00011:00005",
  "USGS:01206900:00011:00001",
  "USGS:01206900:00011:00006",
  "USGS:01208011:00011:00002",
  "USGS:01208500:00011:00002",
  "USGS:01208500:00011:00003",
  "USGS:01208873:00011:00001",
  "USGS:01208873:00011:00002",
  "USGS:01208925:00011:00001",
  "USGS:01208925:00011:00002",
  "USGS:01208950:00011:00005",
  "USGS:01208950:00011:00006",
  "USGS:01208950:00011:00001",
  "USGS:01208950:00011:00003",
  "USGS:01208990:00011:00001",
  "USGS:01208990:00011:00003",
  "USGS:01209005:00011:00002",
  "USGS:01209005:00011:00001",
  "USGS:01209105:00011:00002",
  "USGS:01209105:00011:00001",
  "USGS:01209500:00011:00002",
  "USGS:01209500:00011:00003",
  "USGS:01209510:00011:00001",
  "USGS:012095493:00011:00001",
  "USGS:012095493:00011:00002",
  "USGS:01209700:00011:00001",
  "USGS:01209700:00011:00002",
  "USGS:01209761:00011:00002",
  "USGS:01209761:00011:00001",
  "USGS:01209788:00011:00001",
  "USGS:01209788:00011:00002",
  "USGS:01209901:00011:00001",
  "USGS:01209901:00011:00002",
  "USGS:01212500:00011:00003",
  "USGS:01212500:00011:00002",
  "USGS:01212500:00011:00001",
  "USGS:02176930:00011:00013",
  "USGS:02176930:00011:00003",
  "USGS:02176930:00011:00002",
  "USGS:02176930:00011:00001",
  "USGS:02178400:00011:00006",
  "USGS:02178400:00011:00002",
  "USGS:02178400:00011:00003",
  "USGS:02181350:00011:00005",
  "USGS:02181350:00011:00004",
  "USGS:02181350:00011:00001",
  "USGS:02181580:00011:00003",
  "USGS:02181580:00011:00002",
  "USGS:02181580:00011:00001",
  "USGS:02188600:00011:00005",
  "USGS:02188600:00011:00002",
  "USGS:02188600:00011:00003",
  "USGS:02191227:00011:00004",
  "USGS:02191227:00011:00001",
  "USGS:02191300:00011:00015",
  "USGS:02191300:00011:00013",
  "USGS:02191300:00011:00003",
  "USGS:15051010:00011:00003",
  "USGS:02191740:00011:00003",
  "USGS:02191740:00011:00002",
  "USGS:02191740:00011:00001",
  "USGS:02191743:00011:00003",
  "USGS:02191743:00011:00002",
  "USGS:02191743:00011:00001",
  "USGS:02192000:00011:00001",
  "USGS:02192000:00011:00002",
  "USGS:15008000:00011:00001",
  "USGS:15008000:00011:00002",
  "USGS:15009000:00011:00003",
  "USGS:15009000:00011:00014",
  "USGS:15009000:00011:00001",
  "USGS:15009000:00011:00002",
  "USGS:15009000:00011:00004",
  "USGS:15019990:00011:00002",
  "USGS:15019990:00011:00004",
  "USGS:15024800:00011:00019",
  "USGS:15024800:00011:00004",
  "USGS:15024800:00011:00002",
  "USGS:15024800:00011:00008",
  "USGS:15041200:00011:00016",
  "USGS:15041200:00011:00018",
  "USGS:15041200:00011:00020",
  "USGS:15041200:00011:00021",
  "USGS:15041200:00011:00017",
  "USGS:15041200:00011:00002",
  "USGS:15041200:00011:00005",
  "USGS:15041200:00011:00007",
  "USGS:15051010:00011:00014",
  "USGS:15051010:00011:00002",
  "USGS:15051010:00011:00005",
  "USGS:15052000:00011:00001",
  "USGS:15052000:00011:00002",
  "USGS:15052500:00011:00014",
  "USGS:15052500:00011:00003",
  "USGS:15052500:00011:00004",
  "USGS:15052500:00011:00005",
  "USGS:15055500:00011:00002",
  "USGS:15055500:00011:00001",
  "USGS:15056210:00011:00001",
  "USGS:15056210:00011:00002",
  "USGS:15056210:00011:00005",
  "USGS:15056210:00011:00003",
  "USGS:15056210:00011:00004",
  "USGS:15056500:00011:00008",
  "USGS:15056500:00011:00002",
  "USGS:15056500:00011:00006",
  "USGS:15056500:00011:00009",
  "USGS:15058700:00011:00001",
  "USGS:15058700:00011:00002",
  "USGS:15058700:00011:00003",
  "USGS:15072000:00011:00004",
  "USGS:15072000:00011:00001",
  "USGS:15072000:00011:00002",
  "USGS:15081497:00011:00006",
  "USGS:15081497:00011:00002",
  "USGS:15081497:00011:00004",
  "USGS:15081497:00011:00008",
  "USGS:410628073413301:00011:00001",
  "USGS:4121480721223:00011:00002",
  "USGS:4121480721223:00011:00003",
  "USGS:4121480721223:00011:00001",
  "USGS:412429073165101:00011:00002",
  "USGS:412825072410501:00011:00001",
  "USGS:412916073121701:00011:00001",
  "USGS:413535072253701:00011:00001",
  "USGS:414741072134501:00011:00001",
  "USGS:414831072173002:00011:00001",
  "USGS:02193500:00011:00014",
  "USGS:02193500:00011:00001",
  "USGS:02193500:00011:00004",
  "USGS:02195320:00011:00006",
  "USGS:02195320:00011:00004",
  "USGS:02195320:00011:00003",
  "USGS:02195520:00011:00001",
  "USGS:021964832:00011:00003",
  "USGS:021964832:00011:00005",
  "USGS:021964832:00011:00001",
  "USGS:02196485:00011:00004",
  "USGS:02196485:00011:00001",
  "USGS:02196835:00011:00003",
  "USGS:02196835:00011:00002",
  "USGS:02196835:00011:00001",
  "USGS:02196838:00011:00007",
  "USGS:02196838:00011:00006",
  "USGS:02196838:00011:00003",
  "USGS:02196838:00011:00004",
  "USGS:02196838:00011:00002",
  "USGS:02196838:00011:00018",
  "USGS:02196838:00011:00001",
  "USGS:02196999:00011:00002",
  "USGS:02196999:00011:00001",
  "USGS:02197000:00011:00001",
  "USGS:02197000:00011:00002",
  "USGS:15302200:00011:00014",
  "USGS:15302200:00011:00016",
  "USGS:15302200:00011:00003",
  "USGS:15302200:00011:00001",
  "USGS:15302200:00011:00013",
  "USGS:15302250:00011:00013",
  "USGS:15302250:00011:00015",
  "USGS:15302250:00011:00003",
  "USGS:15302250:00011:00001",
  "USGS:15302250:00011:00002",
  "USGS:15303900:00011:00002",
  "USGS:15303900:00011:00001",
  "USGS:15304000:00011:00016",
  "USGS:15304000:00011:00002",
  "USGS:15304000:00011:00003",
  "USGS:15304010:00011:00001",
  "USGS:15304010:00011:00002",
  "USGS:15320100:00011:00002",
  "USGS:15320100:00011:00001",
  "USGS:15348000:00011:00017",
  "USGS:15348000:00011:00001",
  "USGS:15348000:00011:00002",
  "USGS:15356000:00011:00003",
  "USGS:15356000:00011:00006",
  "USGS:15453500:00011:00017",
  "USGS:15453500:00011:00001",
  "USGS:15453500:00011:00003",
  "USGS:15457790:00011:00004",
  "USGS:15457790:00011:00001",
  "USGS:15457790:00011:00002",
  "USGS:15457800:00011:00001",
  "USGS:15457800:00011:00004",
  "USGS:15457800:00011:00002",
  "USGS:15457800:00011:00003",
  "USGS:15477740:00011:00015",
  "USGS:15477740:00011:00005",
  "USGS:15477740:00011:00002",
  "USGS:15477740:00011:00001",
  "USGS:15478038:00011:00002",
  "USGS:15478038:00011:00004",
  "USGS:15478038:00011:00014",
  "USGS:15478038:00011:00016",
  "USGS:15478038:00011:00020",
  "USGS:15478038:00011:00025",
  "USGS:15478038:00011:00019",
  "USGS:15478038:00011:00001",
  "USGS:15478038:00011:00023",
  "USGS:15478040:00011:00015",
  "USGS:15478040:00011:00016",
  "USGS:15478040:00011:00001",
  "USGS:15478040:00011:00002",
  "USGS:15484000:00011:00019",
  "USGS:15484000:00011:00015",
  "USGS:15484000:00011:00001",
  "USGS:15484000:00011:00002",
  "USGS:15485500:00011:00001",
  "USGS:15485500:00011:00002",
  "USGS:15493000:00011:00021",
  "USGS:15493000:00011:00022",
  "USGS:15493000:00011:00009",
  "USGS:15493000:00011:00001",
  "USGS:15493000:00011:00007",
  "USGS:15493000:00011:00023",
  "USGS:15502000:00011:00012",
  "USGS:15502000:00011:00014",
  "USGS:15502000:00011:00001",
  "USGS:15511000:00011:00020",
  "USGS:15511000:00011:00019",
  "USGS:15511000:00011:00002",
  "USGS:15511000:00011:00006",
  "USGS:15514000:00011:00002",
  "USGS:15514000:00011:00003",
  "USGS:15515060:00011:00003",
  "USGS:15515060:00011:00005",
  "USGS:15515060:00011:00001",
  "USGS:15515060:00011:00002",
  "USGS:15515500:00011:00001",
  "USGS:15515500:00011:00002",
  "USGS:15515500:00011:00003",
  "USGS:15519100:00011:00003",
  "USGS:15519100:00011:00014",
  "USGS:15519100:00011:00001",
  "USGS:15519100:00011:00002",
  "USGS:15519150:00011:00001",
  "USGS:15519150:00011:00002",
  "USGS:15564879:00011:00004",
  "USGS:15564879:00011:00002",
  "USGS:15564879:00011:00003",
  "USGS:15565447:00011:00001",
  "USGS:15565447:00011:00015",
  "USGS:15565447:00011:00002",
  "USGS:15565447:00011:00003",
  "USGS:15580095:00011:00003",
  "USGS:15580095:00011:00004",
  "USGS:15580095:00011:00002",
  "USGS:15580095:00011:00001",
  "USGS:15742980:00011:00002",
  "USGS:15743850:00011:00005",
  "USGS:15743850:00011:00017",
  "USGS:15743850:00011:00002",
  "USGS:15743850:00011:00001",
  "USGS:15744500:00011:00005",
  "USGS:15744500:00011:00006",
  "USGS:15747000:00011:00014",
  "USGS:15747000:00011:00015",
  "USGS:15747000:00011:00004",
  "USGS:15747000:00011:00002",
  "USGS:15803000:00011:00003",
  "USGS:15803000:00011:00004",
  "USGS:15803000:00011:00016",
  "USGS:15803000:00011:00001",
  "USGS:15803000:00011:00002",
  "USGS:15803000:00011:00014",
  "USGS:15820000:00011:00002",
  "USGS:15820000:00011:00014",
  "USGS:15875000:00011:00014",
  "USGS:15875000:00011:00004",
  "USGS:15875000:00011:00001",
  "USGS:15875000:00011:00015",
  "USGS:15875000:00011:00017",
  "USGS:15896000:00011:00001",
  "USGS:15896000:00011:00002",
  "USGS:15896000:00011:00003",
  "USGS:15905100:00011:00004",
  "USGS:15905100:00011:00003",
  "USGS:15905100:00011:00001",
  "USGS:15905100:00011:00002",
  "USGS:15908000:00011:00018",
  "USGS:15908000:00011:00015",
  "USGS:15908000:00011:00014",
  "USGS:15908000:00011:00001",
  "USGS:15908000:00011:00003",
  "USGS:15980000:00011:00004",
  "USGS:15980000:00011:00005",
  "USGS:15980000:00011:00001",
  "USGS:15980000:00011:00002",
  "USGS:16010000:00011:00001",
  "USGS:16010000:00011:00002",
  "USGS:611725149335401:00011:00001",
  "USGS:644528147131202:00011:00001",
  "USGS:644528147131202:00011:00003",
  "USGS:02197020:00011:00003",
  "USGS:02197020:00011:00002",
  "USGS:02197020:00011:00001",
  "USGS:021973269:00011:00003",
  "USGS:021973269:00011:00002",
  "USGS:021973269:00011:00001",
  "USGS:02197500:00011:00001",
  "USGS:02197500:00011:00003",
  "USGS:02197500:00011:00002",
  "USGS:02197598:00011:00002"